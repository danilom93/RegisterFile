
library IEEE;

use IEEE.std_logic_1164.all;

package 
   CONV_PACK_windowedRegisterFile_size_word32_m_global5_n_in_out_local2_f_windows4_size_ext_addr4 
   is

-- define attributes
attribute ENUM_ENCODING : STRING;

end 
   CONV_PACK_windowedRegisterFile_size_word32_m_global5_n_in_out_local2_f_windows4_size_ext_addr4;

library IEEE;

use IEEE.std_logic_1164.all;

use 
   work.CONV_PACK_windowedRegisterFile_size_word32_m_global5_n_in_out_local2_f_windows4_size_ext_addr4.all;

entity register_file_nBitsData32_nBitsAddr5 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end register_file_nBitsData32_nBitsAddr5;

architecture SYN_A of register_file_nBitsData32_nBitsAddr5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
      n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, 
      n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, 
      n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, 
      n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, 
      n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, 
      n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, 
      n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, 
      n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, 
      n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, 
      n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, 
      n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, 
      n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2983, n2984, 
      n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, 
      n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, 
      n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, 
      n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, 
      n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, 
      n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, 
      n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, 
      n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, 
      n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, 
      n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, 
      n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, 
      n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, 
      n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, 
      n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, 
      n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, 
      n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, 
      n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, 
      n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, 
      n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, 
      n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, 
      n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, 
      n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, 
      n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, 
      n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, 
      n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, 
      n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, 
      n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, 
      n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, 
      n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, 
      n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, 
      n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, 
      n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, 
      n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, 
      n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, 
      n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, 
      n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, 
      n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, 
      n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, 
      n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, 
      n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, 
      n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, 
      n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, 
      n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, 
      n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, 
      n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, 
      n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, 
      n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, 
      n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, 
      n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, 
      n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, 
      n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, 
      n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, 
      n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, 
      n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, 
      n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, 
      n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, 
      n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, 
      n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, 
      n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, 
      n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, 
      n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, 
      n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, 
      n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, 
      n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, 
      n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, 
      n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, 
      n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, 
      n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, 
      n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, 
      n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, 
      n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, 
      n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, 
      n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, 
      n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, 
      n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, 
      n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, 
      n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, 
      n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, 
      n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, 
      n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, 
      n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, 
      n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, 
      n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, 
      n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, 
      n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, 
      n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, 
      n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, 
      n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, 
      n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, 
      n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, 
      n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, 
      n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, 
      n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, 
      n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, 
      n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, 
      n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, 
      n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, 
      n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, 
      n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, 
      n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, 
      n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, 
      n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, 
      n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, 
      n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, 
      n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, 
      n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, 
      n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, 
      n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, 
      n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, 
      n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, 
      n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, 
      n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, 
      n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, 
      n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, 
      n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n1,
      n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, 
      n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61
      , n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, 
      n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90
      , n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, 
      n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, 
      n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
      n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
      n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, 
      n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, 
      n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, 
      n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, 
      n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, 
      n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, 
      n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, 
      n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, 
      n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, 
      n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, 
      n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, 
      n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, 
      n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, 
      n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, 
      n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, 
      n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, 
      n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, 
      n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, 
      n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, 
      n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, 
      n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, 
      n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, 
      n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, 
      n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, 
      n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, 
      n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, 
      n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, 
      n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, 
      n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, 
      n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, 
      n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, 
      n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, 
      n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, 
      n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, 
      n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, 
      n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, 
      n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, 
      n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, 
      n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, 
      n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, 
      n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, 
      n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, 
      n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, 
      n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, 
      n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, 
      n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, 
      n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, 
      n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, 
      n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, 
      n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, 
      n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, 
      n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, 
      n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, 
      n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, 
      n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, 
      n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, 
      n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, 
      n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, 
      n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, 
      n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, 
      n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, 
      n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, 
      n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, 
      n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, 
      n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, 
      n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
      n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, 
      n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, 
      n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, 
      n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, 
      n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, 
      n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, 
      n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, 
      n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, 
      n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, 
      n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, 
      n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, 
      n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, 
      n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, 
      n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, 
      n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, 
      n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, 
      n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, 
      n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, 
      n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, 
      n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, 
      n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, 
      n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, 
      n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, 
      n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, 
      n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, 
      n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, 
      n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, 
      n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, 
      n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, 
      n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, 
      n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, 
      n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, 
      n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, 
      n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, 
      n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, 
      n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, 
      n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, 
      n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, 
      n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, 
      n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, 
      n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, 
      n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, 
      n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, 
      n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, 
      n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, 
      n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, 
      n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, 
      n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, 
      n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, 
      n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, 
      n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, 
      n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, 
      n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, 
      n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, 
      n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, 
      n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, 
      n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, 
      n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, 
      n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, 
      n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, 
      n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, 
      n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, 
      n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, 
      n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, 
      n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, 
      n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, 
      n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, 
      n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, 
      n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, 
      n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, 
      n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, 
      n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, 
      n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, 
      n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, 
      n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, 
      n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, 
      n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, 
      n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, 
      n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, 
      n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, 
      n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, 
      n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, 
      n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, 
      n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, 
      n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, 
      n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, 
      n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, 
      n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, 
      n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, 
      n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, 
      n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, 
      n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, 
      n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, 
      n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, 
      n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, 
      n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, 
      n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, 
      n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, 
      n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, 
      n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, 
      n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, 
      n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, 
      n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, 
      n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, 
      n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, 
      n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, 
      n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, 
      n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, 
      n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, 
      n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, 
      n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, 
      n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, 
      n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, 
      n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, 
      n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, 
      n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, 
      n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, 
      n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, 
      n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, 
      n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, 
      n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, 
      n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, 
      n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, 
      n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, 
      n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, 
      n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, 
      n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, 
      n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, 
      n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, 
      n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, 
      n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, 
      n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, 
      n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, 
      n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, 
      n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, 
      n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, 
      n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, 
      n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, 
      n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, 
      n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, 
      n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, 
      n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, 
      n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, 
      n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, 
      n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, 
      n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, 
      n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, 
      n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, 
      n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, 
      n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, 
      n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, 
      n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, 
      n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, 
      n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, 
      n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, 
      n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, 
      n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, 
      n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, 
      n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, 
      n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, 
      n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, 
      n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, 
      n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, 
      n2723, n2724, n2725, n2726, n2855, n2856, n2857, n2858, n2859, n2860, 
      n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, 
      n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, 
      n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, 
      n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, 
      n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, 
      n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, 
      n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, 
      n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, 
      n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, 
      n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, 
      n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, 
      n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, 
      n2981, n2982, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, 
      n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, 
      n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, 
      n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, 
      n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, 
      n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, 
      n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, 
      n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, 
      n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, 
      n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, 
      n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, 
      n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, 
      n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, 
      n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, 
      n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, 
      n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, 
      n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, 
      n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, 
      n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, 
      n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, 
      n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, 
      n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, 
      n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, 
      n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, 
      n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, 
      n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, 
      n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, 
      n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, 
      n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, 
      n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, 
      n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, 
      n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, 
      n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, 
      n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, 
      n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, 
      n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, 
      n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, 
      n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, 
      n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, 
      n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, 
      n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, 
      n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, 
      n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, 
      n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, 
      n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, 
      n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, 
      n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, 
      n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, 
      n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, 
      n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, 
      n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, 
      n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, 
      n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, 
      n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, 
      n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, 
      n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, 
      n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, 
      n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, 
      n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, 
      n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, 
      n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, 
      n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, 
      n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, 
      n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, 
      n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, 
      n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, 
      n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, 
      n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, 
      n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, 
      n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, 
      n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, 
      n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, 
      n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, 
      n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, 
      n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, 
      n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, 
      n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, 
      n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, 
      n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, 
      n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, 
      n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, 
      n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, 
      n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, 
      n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, 
      n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, 
      n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, 
      n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, 
      n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, 
      n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, 
      n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, 
      n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, 
      n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, 
      n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, 
      n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, 
      n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, 
      n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, 
      n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, 
      n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, 
      n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, 
      n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, 
      n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, 
      n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, 
      n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, 
      n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, 
      n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, 
      n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, 
      n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, 
      n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, 
      n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, 
      n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, 
      n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, 
      n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, 
      n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, 
      n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, 
      n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, 
      n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, 
      n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, 
      n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, 
      n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, 
      n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, 
      n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, 
      n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, 
      n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, 
      n5363 : std_logic;

begin
   
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n4102, CK => CLK, Q => n749,
                           QN => n5363);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n4101, CK => CLK, Q => n752,
                           QN => n5362);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n4100, CK => CLK, Q => n754,
                           QN => n5361);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n4099, CK => CLK, Q => n756,
                           QN => n5360);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n4098, CK => CLK, Q => n758,
                           QN => n5359);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n4097, CK => CLK, Q => n760,
                           QN => n5358);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n4096, CK => CLK, Q => n762,
                           QN => n5357);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n4095, CK => CLK, Q => n764,
                           QN => n5356);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n4094, CK => CLK, Q => n766,
                           QN => n5355);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n4093, CK => CLK, Q => n768,
                           QN => n5354);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n4092, CK => CLK, Q => n770,
                           QN => n5353);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n4091, CK => CLK, Q => n772,
                           QN => n5352);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n4090, CK => CLK, Q => n774,
                           QN => n5351);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n4089, CK => CLK, Q => n776,
                           QN => n5350);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n4088, CK => CLK, Q => n778,
                           QN => n5349);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n4087, CK => CLK, Q => n780,
                           QN => n5348);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n4086, CK => CLK, Q => n782,
                           QN => n5347);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n4085, CK => CLK, Q => n784,
                           QN => n5346);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n4084, CK => CLK, Q => n786,
                           QN => n5345);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n4083, CK => CLK, Q => n788,
                           QN => n5344);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n4082, CK => CLK, Q => n790,
                           QN => n5343);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n4081, CK => CLK, Q => n792,
                           QN => n5342);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n4080, CK => CLK, Q => n794, 
                           QN => n5341);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n4079, CK => CLK, Q => n796, 
                           QN => n5340);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n4078, CK => CLK, Q => n798, 
                           QN => n5339);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n4077, CK => CLK, Q => n800, 
                           QN => n5338);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n4076, CK => CLK, Q => n802, 
                           QN => n5337);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n4075, CK => CLK, Q => n804, 
                           QN => n5336);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n4074, CK => CLK, Q => n806, 
                           QN => n5335);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n4073, CK => CLK, Q => n808, 
                           QN => n5334);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n4072, CK => CLK, Q => n810, 
                           QN => n5333);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n4071, CK => CLK, Q => n812, 
                           QN => n5332);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n4070, CK => CLK, Q => n816,
                           QN => n5331);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n4069, CK => CLK, Q => n818,
                           QN => n5330);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n4068, CK => CLK, Q => n819,
                           QN => n5329);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n4067, CK => CLK, Q => n820,
                           QN => n5328);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n4066, CK => CLK, Q => n821,
                           QN => n5327);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n4065, CK => CLK, Q => n822,
                           QN => n5326);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n4064, CK => CLK, Q => n823,
                           QN => n5325);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n4063, CK => CLK, Q => n824,
                           QN => n5324);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n4062, CK => CLK, Q => n825,
                           QN => n5323);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n4061, CK => CLK, Q => n826,
                           QN => n5322);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n4060, CK => CLK, Q => n827,
                           QN => n5321);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n4059, CK => CLK, Q => n828,
                           QN => n5320);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n4058, CK => CLK, Q => n829,
                           QN => n5319);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n4057, CK => CLK, Q => n830,
                           QN => n5318);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n4056, CK => CLK, Q => n831,
                           QN => n5317);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n4055, CK => CLK, Q => n832,
                           QN => n5316);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n4054, CK => CLK, Q => n833,
                           QN => n5315);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n4053, CK => CLK, Q => n834,
                           QN => n5314);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n4052, CK => CLK, Q => n835,
                           QN => n5313);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n4051, CK => CLK, Q => n836,
                           QN => n5312);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n4050, CK => CLK, Q => n837,
                           QN => n5311);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n4049, CK => CLK, Q => n838,
                           QN => n5310);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n4048, CK => CLK, Q => n839, 
                           QN => n5309);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n4047, CK => CLK, Q => n840, 
                           QN => n5308);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n4046, CK => CLK, Q => n841, 
                           QN => n5307);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n4045, CK => CLK, Q => n842, 
                           QN => n5306);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n4044, CK => CLK, Q => n843, 
                           QN => n5305);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n4043, CK => CLK, Q => n844, 
                           QN => n5304);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n4042, CK => CLK, Q => n845, 
                           QN => n5303);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n4041, CK => CLK, Q => n846, 
                           QN => n5302);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n4040, CK => CLK, Q => n847, 
                           QN => n5301);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n4039, CK => CLK, Q => n848, 
                           QN => n5300);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n3974, CK => CLK, Q => n857,
                           QN => n5235);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n3973, CK => CLK, Q => n859,
                           QN => n5234);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n3972, CK => CLK, Q => n860,
                           QN => n5233);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n3971, CK => CLK, Q => n861,
                           QN => n5232);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n3970, CK => CLK, Q => n862,
                           QN => n5231);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n3969, CK => CLK, Q => n863,
                           QN => n5230);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n3968, CK => CLK, Q => n864,
                           QN => n5229);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n3967, CK => CLK, Q => n865,
                           QN => n5228);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n3966, CK => CLK, Q => n866,
                           QN => n5227);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n3965, CK => CLK, Q => n867,
                           QN => n5226);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n3964, CK => CLK, Q => n868,
                           QN => n5225);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n3963, CK => CLK, Q => n869,
                           QN => n5224);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n3962, CK => CLK, Q => n870,
                           QN => n5223);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n3961, CK => CLK, Q => n871,
                           QN => n5222);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n3960, CK => CLK, Q => n872,
                           QN => n5221);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n3959, CK => CLK, Q => n873,
                           QN => n5220);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n3958, CK => CLK, Q => n874,
                           QN => n5219);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n3957, CK => CLK, Q => n875,
                           QN => n5218);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n3956, CK => CLK, Q => n876,
                           QN => n5217);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n3955, CK => CLK, Q => n877,
                           QN => n5216);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n3954, CK => CLK, Q => n878,
                           QN => n5215);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n3953, CK => CLK, Q => n879,
                           QN => n5214);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n3952, CK => CLK, Q => n880, 
                           QN => n5213);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n3951, CK => CLK, Q => n881, 
                           QN => n5212);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n3950, CK => CLK, Q => n882, 
                           QN => n5211);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n3949, CK => CLK, Q => n883, 
                           QN => n5210);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n3948, CK => CLK, Q => n884, 
                           QN => n5209);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n3947, CK => CLK, Q => n885, 
                           QN => n5208);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n3946, CK => CLK, Q => n886, 
                           QN => n5207);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n3945, CK => CLK, Q => n887, 
                           QN => n5206);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n3944, CK => CLK, Q => n888, 
                           QN => n5205);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n3943, CK => CLK, Q => n889, 
                           QN => n5204);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n3942, CK => CLK, Q => n891,
                           QN => n5203);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n3941, CK => CLK, Q => n893,
                           QN => n5202);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n3940, CK => CLK, Q => n894,
                           QN => n5201);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n3939, CK => CLK, Q => n895,
                           QN => n5200);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n3938, CK => CLK, Q => n896,
                           QN => n5199);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n3937, CK => CLK, Q => n897,
                           QN => n5198);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n3936, CK => CLK, Q => n898,
                           QN => n5197);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n3935, CK => CLK, Q => n899,
                           QN => n5196);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n3934, CK => CLK, Q => n900,
                           QN => n5195);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n3933, CK => CLK, Q => n901,
                           QN => n5194);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n3932, CK => CLK, Q => n902,
                           QN => n5193);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n3931, CK => CLK, Q => n903,
                           QN => n5192);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n3930, CK => CLK, Q => n904,
                           QN => n5191);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n3929, CK => CLK, Q => n905,
                           QN => n5190);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n3928, CK => CLK, Q => n906,
                           QN => n5189);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n3927, CK => CLK, Q => n907,
                           QN => n5188);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n3926, CK => CLK, Q => n908,
                           QN => n5187);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n3925, CK => CLK, Q => n909,
                           QN => n5186);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n3924, CK => CLK, Q => n910,
                           QN => n5185);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n3923, CK => CLK, Q => n911,
                           QN => n5184);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n3922, CK => CLK, Q => n912,
                           QN => n5183);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n3921, CK => CLK, Q => n913,
                           QN => n5182);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n3920, CK => CLK, Q => n914, 
                           QN => n5181);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n3919, CK => CLK, Q => n915, 
                           QN => n5180);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n3918, CK => CLK, Q => n916, 
                           QN => n5179);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n3917, CK => CLK, Q => n917, 
                           QN => n5178);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n3916, CK => CLK, Q => n918, 
                           QN => n5177);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n3915, CK => CLK, Q => n919, 
                           QN => n5176);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n3914, CK => CLK, Q => n920, 
                           QN => n5175);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n3913, CK => CLK, Q => n921, 
                           QN => n5174);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n3912, CK => CLK, Q => n922, 
                           QN => n5173);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n3911, CK => CLK, Q => n923, 
                           QN => n5172);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n3846, CK => CLK, Q => n926,
                           QN => n5107);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n3845, CK => CLK, Q => n928,
                           QN => n5106);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n3844, CK => CLK, Q => n929,
                           QN => n5105);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n3843, CK => CLK, Q => n930,
                           QN => n5104);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n3842, CK => CLK, Q => n931,
                           QN => n5103);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n3841, CK => CLK, Q => n932,
                           QN => n5102);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n3840, CK => CLK, Q => n933,
                           QN => n5101);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n3839, CK => CLK, Q => n934,
                           QN => n5100);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n3838, CK => CLK, Q => n935,
                           QN => n5099);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n3837, CK => CLK, Q => n936,
                           QN => n5098);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n3836, CK => CLK, Q => n937,
                           QN => n5097);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n3835, CK => CLK, Q => n938,
                           QN => n5096);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n3834, CK => CLK, Q => n939,
                           QN => n5095);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n3833, CK => CLK, Q => n940,
                           QN => n5094);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n3832, CK => CLK, Q => n941,
                           QN => n5093);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n3831, CK => CLK, Q => n942,
                           QN => n5092);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n3830, CK => CLK, Q => n943,
                           QN => n5091);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n3829, CK => CLK, Q => n944,
                           QN => n5090);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n3828, CK => CLK, Q => n945,
                           QN => n5089);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n3827, CK => CLK, Q => n946,
                           QN => n5088);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n3826, CK => CLK, Q => n947,
                           QN => n5087);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n3825, CK => CLK, Q => n948,
                           QN => n5086);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n3824, CK => CLK, Q => n949, 
                           QN => n5085);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n3823, CK => CLK, Q => n950, 
                           QN => n5084);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n3822, CK => CLK, Q => n951, 
                           QN => n5083);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n3821, CK => CLK, Q => n952, 
                           QN => n5082);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n3820, CK => CLK, Q => n953, 
                           QN => n5081);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n3819, CK => CLK, Q => n954, 
                           QN => n5080);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n3818, CK => CLK, Q => n955, 
                           QN => n5079);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n3817, CK => CLK, Q => n956, 
                           QN => n5078);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n3816, CK => CLK, Q => n957, 
                           QN => n5077);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n3815, CK => CLK, Q => n958, 
                           QN => n5076);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n3814, CK => CLK, Q => n960,
                           QN => n5075);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n3813, CK => CLK, Q => n962,
                           QN => n5074);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n3812, CK => CLK, Q => n963,
                           QN => n5073);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n3811, CK => CLK, Q => n964,
                           QN => n5072);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n3810, CK => CLK, Q => n965,
                           QN => n5071);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n3809, CK => CLK, Q => n966,
                           QN => n5070);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n3808, CK => CLK, Q => n967,
                           QN => n5069);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n3807, CK => CLK, Q => n968,
                           QN => n5068);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n3806, CK => CLK, Q => n969,
                           QN => n5067);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n3805, CK => CLK, Q => n970,
                           QN => n5066);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n3804, CK => CLK, Q => n971,
                           QN => n5065);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n3803, CK => CLK, Q => n972,
                           QN => n5064);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n3802, CK => CLK, Q => n973,
                           QN => n5063);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n3801, CK => CLK, Q => n974,
                           QN => n5062);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n3800, CK => CLK, Q => n975,
                           QN => n5061);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n3799, CK => CLK, Q => n976,
                           QN => n5060);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n3798, CK => CLK, Q => n977,
                           QN => n5059);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n3797, CK => CLK, Q => n978,
                           QN => n5058);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n3796, CK => CLK, Q => n979,
                           QN => n5057);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n3795, CK => CLK, Q => n980,
                           QN => n5056);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n3794, CK => CLK, Q => n981,
                           QN => n5055);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n3793, CK => CLK, Q => n982,
                           QN => n5054);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n3792, CK => CLK, Q => n983, 
                           QN => n5053);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n3791, CK => CLK, Q => n984, 
                           QN => n5052);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n3790, CK => CLK, Q => n985, 
                           QN => n5051);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n3789, CK => CLK, Q => n986, 
                           QN => n5050);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n3788, CK => CLK, Q => n987, 
                           QN => n5049);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n3787, CK => CLK, Q => n988, 
                           QN => n5048);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n3786, CK => CLK, Q => n989, 
                           QN => n5047);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n3785, CK => CLK, Q => n990, 
                           QN => n5046);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n3784, CK => CLK, Q => n991, 
                           QN => n5045);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n3783, CK => CLK, Q => n992, 
                           QN => n5044);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n3718, CK => CLK, Q => n995
                           , QN => n4979);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n3717, CK => CLK, Q => n997
                           , QN => n4978);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n3716, CK => CLK, Q => n998
                           , QN => n4977);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n3715, CK => CLK, Q => n999
                           , QN => n4976);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n3714, CK => CLK, Q => 
                           n1000, QN => n4975);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n3713, CK => CLK, Q => 
                           n1001, QN => n4974);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n3712, CK => CLK, Q => 
                           n1002, QN => n4973);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n3711, CK => CLK, Q => 
                           n1003, QN => n4972);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n3710, CK => CLK, Q => 
                           n1004, QN => n4971);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n3709, CK => CLK, Q => 
                           n1005, QN => n4970);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n3708, CK => CLK, Q => 
                           n1006, QN => n4969);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n3707, CK => CLK, Q => 
                           n1007, QN => n4968);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n3706, CK => CLK, Q => 
                           n1008, QN => n4967);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n3705, CK => CLK, Q => 
                           n1009, QN => n4966);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n3704, CK => CLK, Q => 
                           n1010, QN => n4965);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n3703, CK => CLK, Q => 
                           n1011, QN => n4964);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n3702, CK => CLK, Q => 
                           n1012, QN => n4963);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n3701, CK => CLK, Q => 
                           n1013, QN => n4962);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n3700, CK => CLK, Q => 
                           n1014, QN => n4961);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n3699, CK => CLK, Q => 
                           n1015, QN => n4960);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n3698, CK => CLK, Q => 
                           n1016, QN => n4959);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n3697, CK => CLK, Q => 
                           n1017, QN => n4958);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n3696, CK => CLK, Q => n1018
                           , QN => n4957);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n3695, CK => CLK, Q => n1019
                           , QN => n4956);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n3694, CK => CLK, Q => n1020
                           , QN => n4955);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n3693, CK => CLK, Q => n1021
                           , QN => n4954);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n3692, CK => CLK, Q => n1022
                           , QN => n4953);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n3691, CK => CLK, Q => n1023
                           , QN => n4952);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n3690, CK => CLK, Q => n1024
                           , QN => n4951);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n3689, CK => CLK, Q => n1025
                           , QN => n4950);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n3688, CK => CLK, Q => n1026
                           , QN => n4949);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n3687, CK => CLK, Q => n1027
                           , QN => n4948);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n3686, CK => CLK, Q => 
                           n1029, QN => n4947);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n3685, CK => CLK, Q => 
                           n1031, QN => n4946);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n3684, CK => CLK, Q => 
                           n1032, QN => n4945);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n3683, CK => CLK, Q => 
                           n1033, QN => n4944);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n3682, CK => CLK, Q => 
                           n1034, QN => n4943);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n3681, CK => CLK, Q => 
                           n1035, QN => n4942);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n3680, CK => CLK, Q => 
                           n1036, QN => n4941);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n3679, CK => CLK, Q => 
                           n1037, QN => n4940);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n3678, CK => CLK, Q => 
                           n1038, QN => n4939);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n3677, CK => CLK, Q => 
                           n1039, QN => n4938);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n3676, CK => CLK, Q => 
                           n1040, QN => n4937);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n3675, CK => CLK, Q => 
                           n1041, QN => n4936);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n3674, CK => CLK, Q => 
                           n1042, QN => n4935);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n3673, CK => CLK, Q => 
                           n1043, QN => n4934);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n3672, CK => CLK, Q => 
                           n1044, QN => n4933);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n3671, CK => CLK, Q => 
                           n1045, QN => n4932);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n3670, CK => CLK, Q => 
                           n1046, QN => n4931);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n3669, CK => CLK, Q => 
                           n1047, QN => n4930);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n3668, CK => CLK, Q => 
                           n1048, QN => n4929);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n3667, CK => CLK, Q => 
                           n1049, QN => n4928);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n3666, CK => CLK, Q => 
                           n1050, QN => n4927);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n3665, CK => CLK, Q => 
                           n1051, QN => n4926);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n3664, CK => CLK, Q => n1052
                           , QN => n4925);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n3663, CK => CLK, Q => n1053
                           , QN => n4924);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n3662, CK => CLK, Q => n1054
                           , QN => n4923);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n3661, CK => CLK, Q => n1055
                           , QN => n4922);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n3660, CK => CLK, Q => n1056
                           , QN => n4921);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n3659, CK => CLK, Q => n1057
                           , QN => n4920);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n3658, CK => CLK, Q => n1058
                           , QN => n4919);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n3657, CK => CLK, Q => n1059
                           , QN => n4918);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n3656, CK => CLK, Q => n1060
                           , QN => n4917);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n3655, CK => CLK, Q => n1061
                           , QN => n4916);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n3590, CK => CLK, Q => 
                           n1065, QN => n4851);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n3589, CK => CLK, Q => 
                           n1067, QN => n4850);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n3588, CK => CLK, Q => 
                           n1068, QN => n4849);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n3587, CK => CLK, Q => 
                           n1069, QN => n4848);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n3586, CK => CLK, Q => 
                           n1070, QN => n4847);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n3585, CK => CLK, Q => 
                           n1071, QN => n4846);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n3584, CK => CLK, Q => 
                           n1072, QN => n4845);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n3583, CK => CLK, Q => 
                           n1073, QN => n4844);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n3582, CK => CLK, Q => 
                           n1074, QN => n4843);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n3581, CK => CLK, Q => 
                           n1075, QN => n4842);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n3580, CK => CLK, Q => 
                           n1076, QN => n4841);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n3579, CK => CLK, Q => 
                           n1077, QN => n4840);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n3578, CK => CLK, Q => 
                           n1078, QN => n4839);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n3577, CK => CLK, Q => 
                           n1079, QN => n4838);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n3576, CK => CLK, Q => 
                           n1080, QN => n4837);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n3575, CK => CLK, Q => 
                           n1081, QN => n4836);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n3574, CK => CLK, Q => 
                           n1082, QN => n4835);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n3573, CK => CLK, Q => 
                           n1083, QN => n4834);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n3572, CK => CLK, Q => 
                           n1084, QN => n4833);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n3571, CK => CLK, Q => 
                           n1085, QN => n4832);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n3570, CK => CLK, Q => 
                           n1086, QN => n4831);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n3569, CK => CLK, Q => 
                           n1087, QN => n4830);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n3568, CK => CLK, Q => n1088
                           , QN => n4829);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n3567, CK => CLK, Q => n1089
                           , QN => n4828);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n3566, CK => CLK, Q => n1090
                           , QN => n4827);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n3565, CK => CLK, Q => n1091
                           , QN => n4826);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n3564, CK => CLK, Q => n1092
                           , QN => n4825);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n3563, CK => CLK, Q => n1093
                           , QN => n4824);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n3562, CK => CLK, Q => n1094
                           , QN => n4823);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n3561, CK => CLK, Q => n1095
                           , QN => n4822);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n3560, CK => CLK, Q => n1096
                           , QN => n4821);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n3559, CK => CLK, Q => n1097
                           , QN => n4820);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n3558, CK => CLK, Q => 
                           n1099, QN => n4819);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n3557, CK => CLK, Q => 
                           n1101, QN => n4818);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n3556, CK => CLK, Q => 
                           n1102, QN => n4817);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n3555, CK => CLK, Q => 
                           n1103, QN => n4816);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n3554, CK => CLK, Q => 
                           n1104, QN => n4815);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n3553, CK => CLK, Q => 
                           n1105, QN => n4814);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n3552, CK => CLK, Q => 
                           n1106, QN => n4813);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n3551, CK => CLK, Q => 
                           n1107, QN => n4812);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n3550, CK => CLK, Q => 
                           n1108, QN => n4811);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n3549, CK => CLK, Q => 
                           n1109, QN => n4810);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n3548, CK => CLK, Q => 
                           n1110, QN => n4809);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n3547, CK => CLK, Q => 
                           n1111, QN => n4808);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n3546, CK => CLK, Q => 
                           n1112, QN => n4807);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n3545, CK => CLK, Q => 
                           n1113, QN => n4806);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n3544, CK => CLK, Q => 
                           n1114, QN => n4805);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n3543, CK => CLK, Q => 
                           n1115, QN => n4804);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n3542, CK => CLK, Q => 
                           n1116, QN => n4803);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n3541, CK => CLK, Q => 
                           n1117, QN => n4802);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n3540, CK => CLK, Q => 
                           n1118, QN => n4801);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n3539, CK => CLK, Q => 
                           n1119, QN => n4800);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n3538, CK => CLK, Q => 
                           n1120, QN => n4799);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n3537, CK => CLK, Q => 
                           n1121, QN => n4798);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n3536, CK => CLK, Q => n1122
                           , QN => n4797);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n3535, CK => CLK, Q => n1123
                           , QN => n4796);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n3534, CK => CLK, Q => n1124
                           , QN => n4795);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n3533, CK => CLK, Q => n1125
                           , QN => n4794);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n3532, CK => CLK, Q => n1126
                           , QN => n4793);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n3531, CK => CLK, Q => n1127
                           , QN => n4792);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n3530, CK => CLK, Q => n1128
                           , QN => n4791);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n3529, CK => CLK, Q => n1129
                           , QN => n4790);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n3528, CK => CLK, Q => n1130
                           , QN => n4789);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n3527, CK => CLK, Q => n1131
                           , QN => n4788);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n3462, CK => CLK, Q => 
                           n1135, QN => n4723);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n3461, CK => CLK, Q => 
                           n1137, QN => n4722);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n3460, CK => CLK, Q => 
                           n1138, QN => n4721);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n3459, CK => CLK, Q => 
                           n1139, QN => n4720);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n3458, CK => CLK, Q => 
                           n1140, QN => n4719);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n3457, CK => CLK, Q => 
                           n1141, QN => n4718);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n3456, CK => CLK, Q => 
                           n1142, QN => n4717);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n3455, CK => CLK, Q => 
                           n1143, QN => n4716);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n3454, CK => CLK, Q => 
                           n1144, QN => n4715);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n3453, CK => CLK, Q => 
                           n1145, QN => n4714);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n3452, CK => CLK, Q => 
                           n1146, QN => n4713);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n3451, CK => CLK, Q => 
                           n1147, QN => n4712);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n3450, CK => CLK, Q => 
                           n1148, QN => n4711);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n3449, CK => CLK, Q => 
                           n1149, QN => n4710);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n3448, CK => CLK, Q => 
                           n1150, QN => n4709);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n3447, CK => CLK, Q => 
                           n1151, QN => n4708);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n3446, CK => CLK, Q => 
                           n1152, QN => n4707);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n3445, CK => CLK, Q => 
                           n1153, QN => n4706);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n3444, CK => CLK, Q => 
                           n1154, QN => n4705);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n3443, CK => CLK, Q => 
                           n1155, QN => n4704);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n3442, CK => CLK, Q => 
                           n1156, QN => n4703);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n3441, CK => CLK, Q => 
                           n1157, QN => n4702);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n3440, CK => CLK, Q => n1158
                           , QN => n4701);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n3439, CK => CLK, Q => n1159
                           , QN => n4700);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n3438, CK => CLK, Q => n1160
                           , QN => n4699);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n3437, CK => CLK, Q => n1161
                           , QN => n4698);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n3436, CK => CLK, Q => n1162
                           , QN => n4697);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n3435, CK => CLK, Q => n1163
                           , QN => n4696);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n3434, CK => CLK, Q => n1164
                           , QN => n4695);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n3433, CK => CLK, Q => n1165
                           , QN => n4694);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n3432, CK => CLK, Q => n1166
                           , QN => n4693);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n3431, CK => CLK, Q => n1167
                           , QN => n4692);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n3430, CK => CLK, Q => 
                           n1169, QN => n4691);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n3429, CK => CLK, Q => 
                           n1171, QN => n4690);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n3428, CK => CLK, Q => 
                           n1172, QN => n4689);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n3427, CK => CLK, Q => 
                           n1173, QN => n4688);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n3426, CK => CLK, Q => 
                           n1174, QN => n4687);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n3425, CK => CLK, Q => 
                           n1175, QN => n4686);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n3424, CK => CLK, Q => 
                           n1176, QN => n4685);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n3423, CK => CLK, Q => 
                           n1177, QN => n4684);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n3422, CK => CLK, Q => 
                           n1178, QN => n4683);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n3421, CK => CLK, Q => 
                           n1179, QN => n4682);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n3420, CK => CLK, Q => 
                           n1180, QN => n4681);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n3419, CK => CLK, Q => 
                           n1181, QN => n4680);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n3418, CK => CLK, Q => 
                           n1182, QN => n4679);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n3417, CK => CLK, Q => 
                           n1183, QN => n4678);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n3416, CK => CLK, Q => 
                           n1184, QN => n4677);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n3415, CK => CLK, Q => 
                           n1185, QN => n4676);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n3414, CK => CLK, Q => 
                           n1186, QN => n4675);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n3413, CK => CLK, Q => 
                           n1187, QN => n4674);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n3412, CK => CLK, Q => 
                           n1188, QN => n4673);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n3411, CK => CLK, Q => 
                           n1189, QN => n4672);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n3410, CK => CLK, Q => 
                           n1190, QN => n4671);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n3409, CK => CLK, Q => 
                           n1191, QN => n4670);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n3408, CK => CLK, Q => n1192
                           , QN => n4669);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n3407, CK => CLK, Q => n1193
                           , QN => n4668);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n3406, CK => CLK, Q => n1194
                           , QN => n4667);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n3405, CK => CLK, Q => n1195
                           , QN => n4666);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n3404, CK => CLK, Q => n1196
                           , QN => n4665);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n3403, CK => CLK, Q => n1197
                           , QN => n4664);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n3402, CK => CLK, Q => n1198
                           , QN => n4663);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n3401, CK => CLK, Q => n1199
                           , QN => n4662);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n3400, CK => CLK, Q => n1200
                           , QN => n4661);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n3399, CK => CLK, Q => n1201
                           , QN => n4660);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n3270, CK => CLK, Q => 
                           n1207, QN => n4531);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n3269, CK => CLK, Q => 
                           n1209, QN => n4530);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n3268, CK => CLK, Q => 
                           n1210, QN => n4529);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n3267, CK => CLK, Q => 
                           n1211, QN => n4528);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n3266, CK => CLK, Q => 
                           n1212, QN => n4527);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n3265, CK => CLK, Q => 
                           n1213, QN => n4526);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n3264, CK => CLK, Q => 
                           n1214, QN => n4525);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n3263, CK => CLK, Q => 
                           n1215, QN => n4524);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n3262, CK => CLK, Q => 
                           n1216, QN => n4523);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n3261, CK => CLK, Q => 
                           n1217, QN => n4522);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n3260, CK => CLK, Q => 
                           n1218, QN => n4521);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n3259, CK => CLK, Q => 
                           n1219, QN => n4520);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n3258, CK => CLK, Q => 
                           n1220, QN => n4519);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n3257, CK => CLK, Q => 
                           n1221, QN => n4518);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n3256, CK => CLK, Q => 
                           n1222, QN => n4517);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n3255, CK => CLK, Q => 
                           n1223, QN => n4516);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n3254, CK => CLK, Q => 
                           n1224, QN => n4515);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n3253, CK => CLK, Q => 
                           n1225, QN => n4514);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n3252, CK => CLK, Q => 
                           n1226, QN => n4513);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n3251, CK => CLK, Q => 
                           n1227, QN => n4512);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n3250, CK => CLK, Q => 
                           n1228, QN => n4511);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n3249, CK => CLK, Q => 
                           n1229, QN => n4510);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n3248, CK => CLK, Q => n1230
                           , QN => n4509);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n3247, CK => CLK, Q => n1231
                           , QN => n4508);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n3246, CK => CLK, Q => n1232
                           , QN => n4507);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n3245, CK => CLK, Q => n1233
                           , QN => n4506);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n3244, CK => CLK, Q => n1234
                           , QN => n4505);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n3243, CK => CLK, Q => n1235
                           , QN => n4504);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n3242, CK => CLK, Q => n1236
                           , QN => n4503);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n3241, CK => CLK, Q => n1237
                           , QN => n4502);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n3240, CK => CLK, Q => n1238
                           , QN => n4501);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n3239, CK => CLK, Q => n1239
                           , QN => n4500);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n3238, CK => CLK, Q => 
                           n1240, QN => n4499);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n3237, CK => CLK, Q => 
                           n1242, QN => n4498);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n3236, CK => CLK, Q => 
                           n1243, QN => n4497);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n3235, CK => CLK, Q => 
                           n1244, QN => n4496);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n3234, CK => CLK, Q => 
                           n1245, QN => n4495);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n3233, CK => CLK, Q => 
                           n1246, QN => n4494);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n3232, CK => CLK, Q => 
                           n1247, QN => n4493);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n3231, CK => CLK, Q => 
                           n1248, QN => n4492);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n3230, CK => CLK, Q => 
                           n1249, QN => n4491);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n3229, CK => CLK, Q => 
                           n1250, QN => n4490);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n3228, CK => CLK, Q => 
                           n1251, QN => n4489);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n3227, CK => CLK, Q => 
                           n1252, QN => n4488);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n3226, CK => CLK, Q => 
                           n1253, QN => n4487);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n3225, CK => CLK, Q => 
                           n1254, QN => n4486);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n3224, CK => CLK, Q => 
                           n1255, QN => n4485);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n3223, CK => CLK, Q => 
                           n1256, QN => n4484);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n3222, CK => CLK, Q => 
                           n1257, QN => n4483);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n3221, CK => CLK, Q => 
                           n1258, QN => n4482);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n3220, CK => CLK, Q => 
                           n1259, QN => n4481);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n3219, CK => CLK, Q => 
                           n1260, QN => n4480);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n3218, CK => CLK, Q => 
                           n1261, QN => n4479);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n3217, CK => CLK, Q => 
                           n1262, QN => n4478);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n3216, CK => CLK, Q => n1263
                           , QN => n4477);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n3215, CK => CLK, Q => n1264
                           , QN => n4476);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n3214, CK => CLK, Q => n1265
                           , QN => n4475);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n3213, CK => CLK, Q => n1266
                           , QN => n4474);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n3212, CK => CLK, Q => n1267
                           , QN => n4473);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n3211, CK => CLK, Q => n1268
                           , QN => n4472);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n3210, CK => CLK, Q => n1269
                           , QN => n4471);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n3209, CK => CLK, Q => n1270
                           , QN => n4470);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n3208, CK => CLK, Q => n1271
                           , QN => n4469);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n3207, CK => CLK, Q => n1272
                           , QN => n4468);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n3142, CK => CLK, Q => 
                           n1278, QN => n4403);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n3141, CK => CLK, Q => 
                           n1280, QN => n4402);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n3140, CK => CLK, Q => 
                           n1281, QN => n4401);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n3139, CK => CLK, Q => 
                           n1282, QN => n4400);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n3138, CK => CLK, Q => 
                           n1283, QN => n4399);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n3137, CK => CLK, Q => 
                           n1284, QN => n4398);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n3136, CK => CLK, Q => 
                           n1285, QN => n4397);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n3135, CK => CLK, Q => 
                           n1286, QN => n4396);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n3134, CK => CLK, Q => 
                           n1287, QN => n4395);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n3133, CK => CLK, Q => 
                           n1288, QN => n4394);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n3132, CK => CLK, Q => 
                           n1289, QN => n4393);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n3131, CK => CLK, Q => 
                           n1290, QN => n4392);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n3130, CK => CLK, Q => 
                           n1291, QN => n4391);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n3129, CK => CLK, Q => 
                           n1292, QN => n4390);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n3128, CK => CLK, Q => 
                           n1293, QN => n4389);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n3127, CK => CLK, Q => 
                           n1294, QN => n4388);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n3126, CK => CLK, Q => 
                           n1295, QN => n4387);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n3125, CK => CLK, Q => 
                           n1296, QN => n4386);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n3124, CK => CLK, Q => 
                           n1297, QN => n4385);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n3123, CK => CLK, Q => 
                           n1298, QN => n4384);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n3122, CK => CLK, Q => 
                           n1299, QN => n4383);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n3121, CK => CLK, Q => 
                           n1300, QN => n4382);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n3120, CK => CLK, Q => n1301
                           , QN => n4381);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n3119, CK => CLK, Q => n1302
                           , QN => n4380);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n3118, CK => CLK, Q => n1303
                           , QN => n4379);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n3117, CK => CLK, Q => n1304
                           , QN => n4378);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n3116, CK => CLK, Q => n1305
                           , QN => n4377);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n3115, CK => CLK, Q => n1306
                           , QN => n4376);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n3114, CK => CLK, Q => n1307
                           , QN => n4375);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n3113, CK => CLK, Q => n1308
                           , QN => n4374);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n3112, CK => CLK, Q => n1309
                           , QN => n4373);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n3111, CK => CLK, Q => n1310
                           , QN => n4372);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n3110, CK => CLK, Q => 
                           n1311, QN => n4371);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n3108, CK => CLK, Q => 
                           n1376, QN => n4370);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n3106, CK => CLK, Q => 
                           n1406, QN => n4369);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n3104, CK => CLK, Q => 
                           n1436, QN => n4368);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n3102, CK => CLK, Q => 
                           n1466, QN => n4367);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n3100, CK => CLK, Q => 
                           n1496, QN => n4366);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n3098, CK => CLK, Q => 
                           n1526, QN => n4365);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n3096, CK => CLK, Q => 
                           n1556, QN => n4364);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n3094, CK => CLK, Q => 
                           n1586, QN => n4363);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n3092, CK => CLK, Q => 
                           n1616, QN => n4362);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n3090, CK => CLK, Q => 
                           n1646, QN => n4361);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n3088, CK => CLK, Q => 
                           n1676, QN => n4360);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n3086, CK => CLK, Q => 
                           n1706, QN => n4359);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n3084, CK => CLK, Q => 
                           n1736, QN => n4358);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n3082, CK => CLK, Q => 
                           n1766, QN => n4357);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n3080, CK => CLK, Q => 
                           n1796, QN => n4356);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n3078, CK => CLK, Q => 
                           n1826, QN => n4355);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n3076, CK => CLK, Q => 
                           n1856, QN => n4354);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n3074, CK => CLK, Q => 
                           n1886, QN => n4353);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n3072, CK => CLK, Q => 
                           n1916, QN => n4352);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n3070, CK => CLK, Q => 
                           n1946, QN => n4351);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n3068, CK => CLK, Q => 
                           n1976, QN => n4350);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n3066, CK => CLK, Q => n2006
                           , QN => n4349);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n3064, CK => CLK, Q => n2036
                           , QN => n4348);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n3062, CK => CLK, Q => n2066
                           , QN => n4347);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n3060, CK => CLK, Q => n2096
                           , QN => n4346);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n3058, CK => CLK, Q => n2126
                           , QN => n4345);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n3056, CK => CLK, Q => n2156
                           , QN => n4344);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n3054, CK => CLK, Q => n2186
                           , QN => n4343);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n3052, CK => CLK, Q => n2216
                           , QN => n4342);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n3050, CK => CLK, Q => n2246
                           , QN => n4341);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n3048, CK => CLK, Q => n2276
                           , QN => n4340);
   OUT1_tri_0_inst : TBUF_X1 port map( A => n2853, EN => n2854, Z => OUT1(0));
   OUT1_tri_1_inst : TBUF_X1 port map( A => n2851, EN => n2852, Z => OUT1(1));
   OUT1_tri_2_inst : TBUF_X1 port map( A => n2849, EN => n2850, Z => OUT1(2));
   OUT1_tri_3_inst : TBUF_X1 port map( A => n2847, EN => n2848, Z => OUT1(3));
   OUT1_tri_4_inst : TBUF_X1 port map( A => n2845, EN => n2846, Z => OUT1(4));
   OUT1_tri_5_inst : TBUF_X1 port map( A => n2843, EN => n2844, Z => OUT1(5));
   OUT1_tri_6_inst : TBUF_X1 port map( A => n2841, EN => n2842, Z => OUT1(6));
   OUT1_tri_7_inst : TBUF_X1 port map( A => n2839, EN => n2840, Z => OUT1(7));
   OUT1_tri_8_inst : TBUF_X1 port map( A => n2837, EN => n2838, Z => OUT1(8));
   OUT1_tri_9_inst : TBUF_X1 port map( A => n2835, EN => n2836, Z => OUT1(9));
   OUT1_tri_10_inst : TBUF_X1 port map( A => n2833, EN => n2834, Z => OUT1(10))
                           ;
   OUT1_tri_11_inst : TBUF_X1 port map( A => n2831, EN => n2832, Z => OUT1(11))
                           ;
   OUT1_tri_12_inst : TBUF_X1 port map( A => n2829, EN => n2830, Z => OUT1(12))
                           ;
   OUT1_tri_13_inst : TBUF_X1 port map( A => n2827, EN => n2828, Z => OUT1(13))
                           ;
   OUT1_tri_14_inst : TBUF_X1 port map( A => n2825, EN => n2826, Z => OUT1(14))
                           ;
   OUT1_tri_15_inst : TBUF_X1 port map( A => n2823, EN => n2824, Z => OUT1(15))
                           ;
   OUT1_tri_16_inst : TBUF_X1 port map( A => n2821, EN => n2822, Z => OUT1(16))
                           ;
   OUT1_tri_17_inst : TBUF_X1 port map( A => n2819, EN => n2820, Z => OUT1(17))
                           ;
   OUT1_tri_18_inst : TBUF_X1 port map( A => n2817, EN => n2818, Z => OUT1(18))
                           ;
   OUT1_tri_19_inst : TBUF_X1 port map( A => n2815, EN => n2816, Z => OUT1(19))
                           ;
   OUT1_tri_20_inst : TBUF_X1 port map( A => n2813, EN => n2814, Z => OUT1(20))
                           ;
   OUT1_tri_21_inst : TBUF_X1 port map( A => n2811, EN => n2812, Z => OUT1(21))
                           ;
   OUT1_tri_22_inst : TBUF_X1 port map( A => n2809, EN => n2810, Z => OUT1(22))
                           ;
   OUT1_tri_23_inst : TBUF_X1 port map( A => n2807, EN => n2808, Z => OUT1(23))
                           ;
   OUT1_tri_24_inst : TBUF_X1 port map( A => n2805, EN => n2806, Z => OUT1(24))
                           ;
   OUT1_tri_25_inst : TBUF_X1 port map( A => n2803, EN => n2804, Z => OUT1(25))
                           ;
   OUT1_tri_26_inst : TBUF_X1 port map( A => n2801, EN => n2802, Z => OUT1(26))
                           ;
   OUT1_tri_27_inst : TBUF_X1 port map( A => n2799, EN => n2800, Z => OUT1(27))
                           ;
   OUT1_tri_28_inst : TBUF_X1 port map( A => n2797, EN => n2798, Z => OUT1(28))
                           ;
   OUT1_tri_29_inst : TBUF_X1 port map( A => n2795, EN => n2796, Z => OUT1(29))
                           ;
   OUT1_tri_30_inst : TBUF_X1 port map( A => n2793, EN => n2794, Z => OUT1(30))
                           ;
   OUT1_tri_31_inst : TBUF_X1 port map( A => n2791, EN => n2792, Z => OUT1(31))
                           ;
   OUT2_tri_0_inst : TBUF_X1 port map( A => n2789, EN => n2790, Z => OUT2(0));
   OUT2_tri_1_inst : TBUF_X1 port map( A => n2787, EN => n2788, Z => OUT2(1));
   OUT2_tri_2_inst : TBUF_X1 port map( A => n2785, EN => n2786, Z => OUT2(2));
   OUT2_tri_3_inst : TBUF_X1 port map( A => n2783, EN => n2784, Z => OUT2(3));
   OUT2_tri_4_inst : TBUF_X1 port map( A => n2781, EN => n2782, Z => OUT2(4));
   OUT2_tri_5_inst : TBUF_X1 port map( A => n2779, EN => n2780, Z => OUT2(5));
   OUT2_tri_6_inst : TBUF_X1 port map( A => n2777, EN => n2778, Z => OUT2(6));
   OUT2_tri_7_inst : TBUF_X1 port map( A => n2775, EN => n2776, Z => OUT2(7));
   OUT2_tri_8_inst : TBUF_X1 port map( A => n2773, EN => n2774, Z => OUT2(8));
   OUT2_tri_9_inst : TBUF_X1 port map( A => n2771, EN => n2772, Z => OUT2(9));
   OUT2_tri_10_inst : TBUF_X1 port map( A => n2769, EN => n2770, Z => OUT2(10))
                           ;
   OUT2_tri_11_inst : TBUF_X1 port map( A => n2767, EN => n2768, Z => OUT2(11))
                           ;
   OUT2_tri_12_inst : TBUF_X1 port map( A => n2765, EN => n2766, Z => OUT2(12))
                           ;
   OUT2_tri_13_inst : TBUF_X1 port map( A => n2763, EN => n2764, Z => OUT2(13))
                           ;
   OUT2_tri_14_inst : TBUF_X1 port map( A => n2761, EN => n2762, Z => OUT2(14))
                           ;
   OUT2_tri_15_inst : TBUF_X1 port map( A => n2759, EN => n2760, Z => OUT2(15))
                           ;
   OUT2_tri_16_inst : TBUF_X1 port map( A => n2757, EN => n2758, Z => OUT2(16))
                           ;
   OUT2_tri_17_inst : TBUF_X1 port map( A => n2755, EN => n2756, Z => OUT2(17))
                           ;
   OUT2_tri_18_inst : TBUF_X1 port map( A => n2753, EN => n2754, Z => OUT2(18))
                           ;
   OUT2_tri_19_inst : TBUF_X1 port map( A => n2751, EN => n2752, Z => OUT2(19))
                           ;
   OUT2_tri_20_inst : TBUF_X1 port map( A => n2749, EN => n2750, Z => OUT2(20))
                           ;
   OUT2_tri_21_inst : TBUF_X1 port map( A => n2747, EN => n2748, Z => OUT2(21))
                           ;
   OUT2_tri_22_inst : TBUF_X1 port map( A => n2745, EN => n2746, Z => OUT2(22))
                           ;
   OUT2_tri_23_inst : TBUF_X1 port map( A => n2743, EN => n2744, Z => OUT2(23))
                           ;
   OUT2_tri_24_inst : TBUF_X1 port map( A => n2741, EN => n2742, Z => OUT2(24))
                           ;
   OUT2_tri_25_inst : TBUF_X1 port map( A => n2739, EN => n2740, Z => OUT2(25))
                           ;
   OUT2_tri_26_inst : TBUF_X1 port map( A => n2737, EN => n2738, Z => OUT2(26))
                           ;
   OUT2_tri_27_inst : TBUF_X1 port map( A => n2735, EN => n2736, Z => OUT2(27))
                           ;
   OUT2_tri_28_inst : TBUF_X1 port map( A => n2733, EN => n2734, Z => OUT2(28))
                           ;
   OUT2_tri_29_inst : TBUF_X1 port map( A => n2731, EN => n2732, Z => OUT2(29))
                           ;
   OUT2_tri_30_inst : TBUF_X1 port map( A => n2729, EN => n2730, Z => OUT2(30))
                           ;
   OUT2_tri_31_inst : TBUF_X1 port map( A => n2727, EN => n2728, Z => OUT2(31))
                           ;
   OUT2_tri_enable_reg_31_inst : DFF_X1 port map( D => n4134, CK => CLK, Q => 
                           n2728, QN => n714);
   OUT2_tri_enable_reg_28_inst : DFF_X1 port map( D => n4131, CK => CLK, Q => 
                           n2734, QN => n718);
   OUT2_tri_enable_reg_27_inst : DFF_X1 port map( D => n4130, CK => CLK, Q => 
                           n2736, QN => n719);
   OUT1_tri_enable_reg_31_inst : DFF_X1 port map( D => n3045, CK => CLK, Q => 
                           n2792, QN => n2383);
   OUT1_tri_enable_reg_30_inst : DFF_X1 port map( D => n3043, CK => CLK, Q => 
                           n2794, QN => n2405);
   OUT1_tri_enable_reg_29_inst : DFF_X1 port map( D => n3041, CK => CLK, Q => 
                           n2796, QN => n2426);
   OUT1_tri_enable_reg_28_inst : DFF_X1 port map( D => n3039, CK => CLK, Q => 
                           n2798, QN => n2447);
   OUT1_tri_enable_reg_27_inst : DFF_X1 port map( D => n3037, CK => CLK, Q => 
                           n2800, QN => n2468);
   OUT1_tri_enable_reg_26_inst : DFF_X1 port map( D => n3035, CK => CLK, Q => 
                           n2802, QN => n2489);
   OUT1_tri_enable_reg_25_inst : DFF_X1 port map( D => n3033, CK => CLK, Q => 
                           n2804, QN => n2510);
   OUT1_tri_enable_reg_24_inst : DFF_X1 port map( D => n3031, CK => CLK, Q => 
                           n2806, QN => n2531);
   OUT2_tri_enable_reg_30_inst : DFF_X1 port map( D => n4133, CK => CLK, Q => 
                           n2730, QN => n716);
   OUT2_tri_enable_reg_29_inst : DFF_X1 port map( D => n4132, CK => CLK, Q => 
                           n2732, QN => n717);
   OUT2_tri_enable_reg_26_inst : DFF_X1 port map( D => n4129, CK => CLK, Q => 
                           n2738, QN => n720);
   OUT2_tri_enable_reg_25_inst : DFF_X1 port map( D => n4128, CK => CLK, Q => 
                           n2740, QN => n721);
   OUT2_tri_enable_reg_24_inst : DFF_X1 port map( D => n4127, CK => CLK, Q => 
                           n2742, QN => n722);
   OUT1_tri_enable_reg_19_inst : DFF_X1 port map( D => n3021, CK => CLK, Q => 
                           n2816, QN => n2636);
   OUT1_tri_enable_reg_17_inst : DFF_X1 port map( D => n3017, CK => CLK, Q => 
                           n2820, QN => n2678);
   OUT1_tri_enable_reg_15_inst : DFF_X1 port map( D => n3013, CK => CLK, Q => 
                           n2824, QN => n2720);
   OUT1_tri_enable_reg_13_inst : DFF_X1 port map( D => n3009, CK => CLK, Q => 
                           n2828, QN => n2890);
   OUT1_tri_enable_reg_11_inst : DFF_X1 port map( D => n3005, CK => CLK, Q => 
                           n2832, QN => n2932);
   OUT1_tri_enable_reg_7_inst : DFF_X1 port map( D => n2997, CK => CLK, Q => 
                           n2840, QN => n4168);
   OUT1_tri_enable_reg_5_inst : DFF_X1 port map( D => n2993, CK => CLK, Q => 
                           n2844, QN => n4210);
   OUT1_tri_enable_reg_3_inst : DFF_X1 port map( D => n2989, CK => CLK, Q => 
                           n2848, QN => n4252);
   OUT1_tri_enable_reg_2_inst : DFF_X1 port map( D => n2987, CK => CLK, Q => 
                           n2850, QN => n4273);
   OUT1_tri_enable_reg_1_inst : DFF_X1 port map( D => n2985, CK => CLK, Q => 
                           n2852, QN => n4294);
   OUT2_tri_enable_reg_23_inst : DFF_X1 port map( D => n4126, CK => CLK, Q => 
                           n2744, QN => n723);
   OUT2_tri_enable_reg_21_inst : DFF_X1 port map( D => n4124, CK => CLK, Q => 
                           n2748, QN => n725);
   OUT2_tri_enable_reg_20_inst : DFF_X1 port map( D => n4123, CK => CLK, Q => 
                           n2750, QN => n726);
   OUT2_tri_enable_reg_19_inst : DFF_X1 port map( D => n4122, CK => CLK, Q => 
                           n2752, QN => n727);
   OUT2_tri_enable_reg_18_inst : DFF_X1 port map( D => n4121, CK => CLK, Q => 
                           n2754, QN => n728);
   OUT2_tri_enable_reg_17_inst : DFF_X1 port map( D => n4120, CK => CLK, Q => 
                           n2756, QN => n729);
   OUT2_tri_enable_reg_16_inst : DFF_X1 port map( D => n4119, CK => CLK, Q => 
                           n2758, QN => n730);
   OUT2_tri_enable_reg_15_inst : DFF_X1 port map( D => n4118, CK => CLK, Q => 
                           n2760, QN => n731);
   OUT2_tri_enable_reg_14_inst : DFF_X1 port map( D => n4117, CK => CLK, Q => 
                           n2762, QN => n732);
   OUT2_tri_enable_reg_13_inst : DFF_X1 port map( D => n4116, CK => CLK, Q => 
                           n2764, QN => n733);
   OUT2_tri_enable_reg_12_inst : DFF_X1 port map( D => n4115, CK => CLK, Q => 
                           n2766, QN => n734);
   OUT2_tri_enable_reg_11_inst : DFF_X1 port map( D => n4114, CK => CLK, Q => 
                           n2768, QN => n735);
   OUT2_tri_enable_reg_10_inst : DFF_X1 port map( D => n4113, CK => CLK, Q => 
                           n2770, QN => n736);
   OUT2_tri_enable_reg_9_inst : DFF_X1 port map( D => n4112, CK => CLK, Q => 
                           n2772, QN => n737);
   OUT2_tri_enable_reg_8_inst : DFF_X1 port map( D => n4111, CK => CLK, Q => 
                           n2774, QN => n738);
   OUT2_tri_enable_reg_7_inst : DFF_X1 port map( D => n4110, CK => CLK, Q => 
                           n2776, QN => n739);
   OUT2_tri_enable_reg_6_inst : DFF_X1 port map( D => n4109, CK => CLK, Q => 
                           n2778, QN => n740);
   OUT2_tri_enable_reg_5_inst : DFF_X1 port map( D => n4108, CK => CLK, Q => 
                           n2780, QN => n741);
   OUT2_tri_enable_reg_4_inst : DFF_X1 port map( D => n4107, CK => CLK, Q => 
                           n2782, QN => n742);
   OUT2_tri_enable_reg_3_inst : DFF_X1 port map( D => n4106, CK => CLK, Q => 
                           n2784, QN => n743);
   OUT2_tri_enable_reg_2_inst : DFF_X1 port map( D => n4105, CK => CLK, Q => 
                           n2786, QN => n744);
   OUT2_tri_enable_reg_1_inst : DFF_X1 port map( D => n4104, CK => CLK, Q => 
                           n2788, QN => n745);
   OUT2_tri_enable_reg_0_inst : DFF_X1 port map( D => n4103, CK => CLK, Q => 
                           n2790, QN => n746);
   OUT1_tri_enable_reg_23_inst : DFF_X1 port map( D => n3029, CK => CLK, Q => 
                           n2808, QN => n2552);
   OUT1_tri_enable_reg_22_inst : DFF_X1 port map( D => n3027, CK => CLK, Q => 
                           n2810, QN => n2573);
   OUT1_tri_enable_reg_21_inst : DFF_X1 port map( D => n3025, CK => CLK, Q => 
                           n2812, QN => n2594);
   OUT1_tri_enable_reg_20_inst : DFF_X1 port map( D => n3023, CK => CLK, Q => 
                           n2814, QN => n2615);
   OUT1_tri_enable_reg_18_inst : DFF_X1 port map( D => n3019, CK => CLK, Q => 
                           n2818, QN => n2657);
   OUT1_tri_enable_reg_16_inst : DFF_X1 port map( D => n3015, CK => CLK, Q => 
                           n2822, QN => n2699);
   OUT1_tri_enable_reg_14_inst : DFF_X1 port map( D => n3011, CK => CLK, Q => 
                           n2826, QN => n2869);
   OUT1_tri_enable_reg_12_inst : DFF_X1 port map( D => n3007, CK => CLK, Q => 
                           n2830, QN => n2911);
   OUT1_tri_enable_reg_10_inst : DFF_X1 port map( D => n3003, CK => CLK, Q => 
                           n2834, QN => n2953);
   OUT1_tri_enable_reg_9_inst : DFF_X1 port map( D => n3001, CK => CLK, Q => 
                           n2836, QN => n2974);
   OUT1_tri_enable_reg_8_inst : DFF_X1 port map( D => n2999, CK => CLK, Q => 
                           n2838, QN => n4147);
   OUT1_tri_enable_reg_6_inst : DFF_X1 port map( D => n2995, CK => CLK, Q => 
                           n2842, QN => n4189);
   OUT1_tri_enable_reg_4_inst : DFF_X1 port map( D => n2991, CK => CLK, Q => 
                           n2846, QN => n4231);
   OUT1_tri_enable_reg_0_inst : DFF_X1 port map( D => n2983, CK => CLK, Q => 
                           n2854, QN => n4339);
   OUT2_tri_enable_reg_22_inst : DFF_X1 port map( D => n4125, CK => CLK, Q => 
                           n2746, QN => n724);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n3174, CK => CLK, Q => 
                           n4435, QN => n1365);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n3173, CK => CLK, Q => 
                           n4434, QN => n1401);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n3172, CK => CLK, Q => 
                           n4433, QN => n1431);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n3171, CK => CLK, Q => 
                           n4432, QN => n1461);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n3170, CK => CLK, Q => 
                           n4431, QN => n1491);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n3169, CK => CLK, Q => 
                           n4430, QN => n1521);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n3168, CK => CLK, Q => 
                           n4429, QN => n1551);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n3167, CK => CLK, Q => 
                           n4428, QN => n1581);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n3206, CK => CLK, Q => 
                           n4467, QN => n1367);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n3205, CK => CLK, Q => 
                           n4466, QN => n1402);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n3204, CK => CLK, Q => 
                           n4465, QN => n1432);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n3203, CK => CLK, Q => 
                           n4464, QN => n1462);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n3202, CK => CLK, Q => 
                           n4463, QN => n1492);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n3201, CK => CLK, Q => 
                           n4462, QN => n1522);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n3200, CK => CLK, Q => 
                           n4461, QN => n1552);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n3199, CK => CLK, Q => 
                           n4460, QN => n1582);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n3334, CK => CLK, Q => 
                           n4595, QN => n256);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n3333, CK => CLK, Q => 
                           n4594, QN => n255);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n3332, CK => CLK, Q => 
                           n4593, QN => n254);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n3331, CK => CLK, Q => 
                           n4592, QN => n253);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n3330, CK => CLK, Q => 
                           n4591, QN => n252);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n3329, CK => CLK, Q => 
                           n4590, QN => n251);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n3328, CK => CLK, Q => 
                           n4589, QN => n250);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n3327, CK => CLK, Q => 
                           n4588, QN => n249);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n3398, CK => CLK, Q => 
                           n4659, QN => n248);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n3397, CK => CLK, Q => 
                           n4658, QN => n247);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n3396, CK => CLK, Q => 
                           n4657, QN => n246);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n3395, CK => CLK, Q => 
                           n4656, QN => n245);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n3394, CK => CLK, Q => 
                           n4655, QN => n244);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n3393, CK => CLK, Q => 
                           n4654, QN => n243);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n3392, CK => CLK, Q => 
                           n4653, QN => n242);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n3391, CK => CLK, Q => 
                           n4652, QN => n241);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n3366, CK => CLK, Q => 
                           n4627, QN => n240);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n3365, CK => CLK, Q => 
                           n4626, QN => n239);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n3364, CK => CLK, Q => 
                           n4625, QN => n238);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n3363, CK => CLK, Q => 
                           n4624, QN => n237);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n3362, CK => CLK, Q => 
                           n4623, QN => n236);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n3361, CK => CLK, Q => 
                           n4622, QN => n235);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n3360, CK => CLK, Q => 
                           n4621, QN => n234);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n3359, CK => CLK, Q => 
                           n4620, QN => n233);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n3494, CK => CLK, Q => 
                           n4755, QN => n1372);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n3493, CK => CLK, Q => 
                           n4754, QN => n1404);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n3492, CK => CLK, Q => 
                           n4753, QN => n1434);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n3491, CK => CLK, Q => 
                           n4752, QN => n1464);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n3490, CK => CLK, Q => 
                           n4751, QN => n1494);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n3489, CK => CLK, Q => 
                           n4750, QN => n1524);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n3488, CK => CLK, Q => 
                           n4749, QN => n1554);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n3487, CK => CLK, Q => 
                           n4748, QN => n1584);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n3302, CK => CLK, Q => 
                           n4563, QN => n232);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n3301, CK => CLK, Q => 
                           n4562, QN => n231);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n3300, CK => CLK, Q => 
                           n4561, QN => n230);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n3299, CK => CLK, Q => 
                           n4560, QN => n229);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n3298, CK => CLK, Q => 
                           n4559, QN => n228);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n3297, CK => CLK, Q => 
                           n4558, QN => n227);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n3296, CK => CLK, Q => 
                           n4557, QN => n226);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n3295, CK => CLK, Q => 
                           n4556, QN => n225);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n3526, CK => CLK, Q => 
                           n4787, QN => n1374);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n3525, CK => CLK, Q => 
                           n4786, QN => n1405);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n3524, CK => CLK, Q => 
                           n4785, QN => n1435);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n3523, CK => CLK, Q => 
                           n4784, QN => n1465);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n3522, CK => CLK, Q => 
                           n4783, QN => n1495);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n3521, CK => CLK, Q => 
                           n4782, QN => n1525);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n3520, CK => CLK, Q => 
                           n4781, QN => n1555);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n3519, CK => CLK, Q => 
                           n4780, QN => n1585);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n3166, CK => CLK, Q => 
                           n4427, QN => n1611);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n3165, CK => CLK, Q => 
                           n4426, QN => n1641);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n3164, CK => CLK, Q => 
                           n4425, QN => n1671);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n3163, CK => CLK, Q => 
                           n4424, QN => n1701);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n3162, CK => CLK, Q => 
                           n4423, QN => n1731);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n3161, CK => CLK, Q => 
                           n4422, QN => n1761);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n3160, CK => CLK, Q => 
                           n4421, QN => n1791);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n3159, CK => CLK, Q => 
                           n4420, QN => n1821);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n3158, CK => CLK, Q => 
                           n4419, QN => n1851);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n3157, CK => CLK, Q => 
                           n4418, QN => n1881);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n3156, CK => CLK, Q => 
                           n4417, QN => n1911);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n3155, CK => CLK, Q => 
                           n4416, QN => n1941);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n3154, CK => CLK, Q => 
                           n4415, QN => n1971);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n3153, CK => CLK, Q => 
                           n4414, QN => n2001);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n3152, CK => CLK, Q => n4413
                           , QN => n2031);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n3151, CK => CLK, Q => n4412
                           , QN => n2061);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n3150, CK => CLK, Q => n4411
                           , QN => n2091);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n3149, CK => CLK, Q => n4410
                           , QN => n2121);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n3148, CK => CLK, Q => n4409
                           , QN => n2151);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n3147, CK => CLK, Q => n4408
                           , QN => n2181);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n3146, CK => CLK, Q => n4407
                           , QN => n2211);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n3145, CK => CLK, Q => n4406
                           , QN => n2241);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n3144, CK => CLK, Q => n4405
                           , QN => n2271);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n3143, CK => CLK, Q => n4404
                           , QN => n2315);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n3198, CK => CLK, Q => 
                           n4459, QN => n1612);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n3197, CK => CLK, Q => 
                           n4458, QN => n1642);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n3196, CK => CLK, Q => 
                           n4457, QN => n1672);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n3195, CK => CLK, Q => 
                           n4456, QN => n1702);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n3194, CK => CLK, Q => 
                           n4455, QN => n1732);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n3193, CK => CLK, Q => 
                           n4454, QN => n1762);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n3192, CK => CLK, Q => 
                           n4453, QN => n1792);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n3191, CK => CLK, Q => 
                           n4452, QN => n1822);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n3190, CK => CLK, Q => 
                           n4451, QN => n1852);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n3189, CK => CLK, Q => 
                           n4450, QN => n1882);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n3188, CK => CLK, Q => 
                           n4449, QN => n1912);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n3187, CK => CLK, Q => 
                           n4448, QN => n1942);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n3186, CK => CLK, Q => 
                           n4447, QN => n1972);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n3185, CK => CLK, Q => 
                           n4446, QN => n2002);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n3184, CK => CLK, Q => n4445
                           , QN => n2032);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n3183, CK => CLK, Q => n4444
                           , QN => n2062);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n3182, CK => CLK, Q => n4443
                           , QN => n2092);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n3181, CK => CLK, Q => n4442
                           , QN => n2122);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n3180, CK => CLK, Q => n4441
                           , QN => n2152);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n3179, CK => CLK, Q => n4440
                           , QN => n2182);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n3178, CK => CLK, Q => n4439
                           , QN => n2212);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n3177, CK => CLK, Q => n4438
                           , QN => n2242);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n3176, CK => CLK, Q => n4437
                           , QN => n2272);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n3175, CK => CLK, Q => n4436
                           , QN => n2316);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n3326, CK => CLK, Q => 
                           n4587, QN => n224);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n3325, CK => CLK, Q => 
                           n4586, QN => n223);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n3324, CK => CLK, Q => 
                           n4585, QN => n222);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n3323, CK => CLK, Q => 
                           n4584, QN => n221);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n3322, CK => CLK, Q => 
                           n4583, QN => n220);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n3321, CK => CLK, Q => 
                           n4582, QN => n219);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n3320, CK => CLK, Q => 
                           n4581, QN => n218);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n3319, CK => CLK, Q => 
                           n4580, QN => n217);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n3318, CK => CLK, Q => 
                           n4579, QN => n216);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n3317, CK => CLK, Q => 
                           n4578, QN => n215);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n3316, CK => CLK, Q => 
                           n4577, QN => n214);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n3315, CK => CLK, Q => 
                           n4576, QN => n213);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n3314, CK => CLK, Q => 
                           n4575, QN => n212);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n3313, CK => CLK, Q => 
                           n4574, QN => n211);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n3312, CK => CLK, Q => n4573
                           , QN => n210);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n3311, CK => CLK, Q => n4572
                           , QN => n209);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n3310, CK => CLK, Q => n4571
                           , QN => n208);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n3309, CK => CLK, Q => n4570
                           , QN => n207);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n3308, CK => CLK, Q => n4569
                           , QN => n206);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n3307, CK => CLK, Q => n4568
                           , QN => n205);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n3306, CK => CLK, Q => n4567
                           , QN => n204);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n3305, CK => CLK, Q => n4566
                           , QN => n203);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n3304, CK => CLK, Q => n4565
                           , QN => n202);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n3303, CK => CLK, Q => n4564
                           , QN => n201);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n3390, CK => CLK, Q => 
                           n4651, QN => n200);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n3389, CK => CLK, Q => 
                           n4650, QN => n199);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n3388, CK => CLK, Q => 
                           n4649, QN => n198);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n3387, CK => CLK, Q => 
                           n4648, QN => n197);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n3386, CK => CLK, Q => 
                           n4647, QN => n196);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n3385, CK => CLK, Q => 
                           n4646, QN => n195);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n3384, CK => CLK, Q => 
                           n4645, QN => n194);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n3383, CK => CLK, Q => 
                           n4644, QN => n193);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n3382, CK => CLK, Q => 
                           n4643, QN => n192);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n3381, CK => CLK, Q => 
                           n4642, QN => n191);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n3380, CK => CLK, Q => 
                           n4641, QN => n190);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n3379, CK => CLK, Q => 
                           n4640, QN => n189);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n3378, CK => CLK, Q => 
                           n4639, QN => n188);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n3377, CK => CLK, Q => 
                           n4638, QN => n187);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n3376, CK => CLK, Q => n4637
                           , QN => n186);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n3375, CK => CLK, Q => n4636
                           , QN => n185);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n3374, CK => CLK, Q => n4635
                           , QN => n184);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n3373, CK => CLK, Q => n4634
                           , QN => n183);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n3372, CK => CLK, Q => n4633
                           , QN => n182);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n3371, CK => CLK, Q => n4632
                           , QN => n181);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n3370, CK => CLK, Q => n4631
                           , QN => n180);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n3369, CK => CLK, Q => n4630
                           , QN => n179);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n3368, CK => CLK, Q => n4629
                           , QN => n178);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n3367, CK => CLK, Q => n4628
                           , QN => n177);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n3358, CK => CLK, Q => 
                           n4619, QN => n176);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n3357, CK => CLK, Q => 
                           n4618, QN => n175);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n3356, CK => CLK, Q => 
                           n4617, QN => n174);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n3355, CK => CLK, Q => 
                           n4616, QN => n173);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n3354, CK => CLK, Q => 
                           n4615, QN => n172);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n3353, CK => CLK, Q => 
                           n4614, QN => n171);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n3352, CK => CLK, Q => 
                           n4613, QN => n170);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n3351, CK => CLK, Q => 
                           n4612, QN => n169);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n3350, CK => CLK, Q => 
                           n4611, QN => n168);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n3349, CK => CLK, Q => 
                           n4610, QN => n167);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n3348, CK => CLK, Q => 
                           n4609, QN => n166);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n3347, CK => CLK, Q => 
                           n4608, QN => n165);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n3346, CK => CLK, Q => 
                           n4607, QN => n164);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n3345, CK => CLK, Q => 
                           n4606, QN => n163);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n3344, CK => CLK, Q => n4605
                           , QN => n162);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n3343, CK => CLK, Q => n4604
                           , QN => n161);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n3342, CK => CLK, Q => n4603
                           , QN => n160);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n3341, CK => CLK, Q => n4602
                           , QN => n159);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n3340, CK => CLK, Q => n4601
                           , QN => n158);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n3339, CK => CLK, Q => n4600
                           , QN => n157);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n3338, CK => CLK, Q => n4599
                           , QN => n156);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n3337, CK => CLK, Q => n4598
                           , QN => n155);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n3336, CK => CLK, Q => n4597
                           , QN => n154);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n3335, CK => CLK, Q => n4596
                           , QN => n153);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n3486, CK => CLK, Q => 
                           n4747, QN => n1614);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n3485, CK => CLK, Q => 
                           n4746, QN => n1644);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n3484, CK => CLK, Q => 
                           n4745, QN => n1674);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n3483, CK => CLK, Q => 
                           n4744, QN => n1704);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n3482, CK => CLK, Q => 
                           n4743, QN => n1734);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n3481, CK => CLK, Q => 
                           n4742, QN => n1764);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n3480, CK => CLK, Q => 
                           n4741, QN => n1794);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n3479, CK => CLK, Q => 
                           n4740, QN => n1824);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n3478, CK => CLK, Q => 
                           n4739, QN => n1854);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n3477, CK => CLK, Q => 
                           n4738, QN => n1884);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n3476, CK => CLK, Q => 
                           n4737, QN => n1914);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n3475, CK => CLK, Q => 
                           n4736, QN => n1944);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n3474, CK => CLK, Q => 
                           n4735, QN => n1974);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n3473, CK => CLK, Q => 
                           n4734, QN => n2004);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n3472, CK => CLK, Q => n4733
                           , QN => n2034);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n3471, CK => CLK, Q => n4732
                           , QN => n2064);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n3470, CK => CLK, Q => n4731
                           , QN => n2094);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n3469, CK => CLK, Q => n4730
                           , QN => n2124);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n3468, CK => CLK, Q => n4729
                           , QN => n2154);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n3467, CK => CLK, Q => n4728
                           , QN => n2184);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n3466, CK => CLK, Q => n4727
                           , QN => n2214);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n3465, CK => CLK, Q => n4726
                           , QN => n2244);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n3464, CK => CLK, Q => n4725
                           , QN => n2274);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n3463, CK => CLK, Q => n4724
                           , QN => n2320);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n3294, CK => CLK, Q => 
                           n4555, QN => n152);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n3293, CK => CLK, Q => 
                           n4554, QN => n151);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n3292, CK => CLK, Q => 
                           n4553, QN => n150);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n3291, CK => CLK, Q => 
                           n4552, QN => n149);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n3290, CK => CLK, Q => 
                           n4551, QN => n148);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n3289, CK => CLK, Q => 
                           n4550, QN => n147);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n3288, CK => CLK, Q => 
                           n4549, QN => n146);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n3287, CK => CLK, Q => 
                           n4548, QN => n145);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n3286, CK => CLK, Q => 
                           n4547, QN => n144);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n3285, CK => CLK, Q => 
                           n4546, QN => n143);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n3284, CK => CLK, Q => 
                           n4545, QN => n142);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n3283, CK => CLK, Q => 
                           n4544, QN => n141);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n3282, CK => CLK, Q => 
                           n4543, QN => n140);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n3281, CK => CLK, Q => 
                           n4542, QN => n139);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n3280, CK => CLK, Q => n4541
                           , QN => n138);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n3279, CK => CLK, Q => n4540
                           , QN => n137);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n3278, CK => CLK, Q => n4539
                           , QN => n136);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n3277, CK => CLK, Q => n4538
                           , QN => n135);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n3276, CK => CLK, Q => n4537
                           , QN => n134);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n3275, CK => CLK, Q => n4536
                           , QN => n133);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n3274, CK => CLK, Q => n4535
                           , QN => n132);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n3273, CK => CLK, Q => n4534
                           , QN => n131);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n3272, CK => CLK, Q => n4533
                           , QN => n130);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n3271, CK => CLK, Q => n4532
                           , QN => n129);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n3518, CK => CLK, Q => 
                           n4779, QN => n1615);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n3517, CK => CLK, Q => 
                           n4778, QN => n1645);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n3516, CK => CLK, Q => 
                           n4777, QN => n1675);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n3515, CK => CLK, Q => 
                           n4776, QN => n1705);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n3514, CK => CLK, Q => 
                           n4775, QN => n1735);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n3513, CK => CLK, Q => 
                           n4774, QN => n1765);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n3512, CK => CLK, Q => 
                           n4773, QN => n1795);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n3511, CK => CLK, Q => 
                           n4772, QN => n1825);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n3510, CK => CLK, Q => 
                           n4771, QN => n1855);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n3509, CK => CLK, Q => 
                           n4770, QN => n1885);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n3508, CK => CLK, Q => 
                           n4769, QN => n1915);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n3507, CK => CLK, Q => 
                           n4768, QN => n1945);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n3506, CK => CLK, Q => 
                           n4767, QN => n1975);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n3505, CK => CLK, Q => 
                           n4766, QN => n2005);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n3504, CK => CLK, Q => n4765
                           , QN => n2035);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n3503, CK => CLK, Q => n4764
                           , QN => n2065);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n3502, CK => CLK, Q => n4763
                           , QN => n2095);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n3501, CK => CLK, Q => n4762
                           , QN => n2125);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n3500, CK => CLK, Q => n4761
                           , QN => n2155);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n3499, CK => CLK, Q => n4760
                           , QN => n2185);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n3498, CK => CLK, Q => n4759
                           , QN => n2215);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n3497, CK => CLK, Q => n4758
                           , QN => n2245);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n3496, CK => CLK, Q => n4757
                           , QN => n2275);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n3495, CK => CLK, Q => n4756
                           , QN => n2321);
   OUT1_reg_31_inst : DFF_X1 port map( D => n3046, CK => CLK, Q => n2791, QN =>
                           n2330);
   OUT1_reg_30_inst : DFF_X1 port map( D => n3044, CK => CLK, Q => n2793, QN =>
                           n2385);
   OUT1_reg_29_inst : DFF_X1 port map( D => n3042, CK => CLK, Q => n2795, QN =>
                           n2406);
   OUT1_reg_28_inst : DFF_X1 port map( D => n3040, CK => CLK, Q => n2797, QN =>
                           n2427);
   OUT1_reg_27_inst : DFF_X1 port map( D => n3038, CK => CLK, Q => n2799, QN =>
                           n2448);
   OUT1_reg_26_inst : DFF_X1 port map( D => n3036, CK => CLK, Q => n2801, QN =>
                           n2469);
   OUT1_reg_25_inst : DFF_X1 port map( D => n3034, CK => CLK, Q => n2803, QN =>
                           n2490);
   OUT1_reg_24_inst : DFF_X1 port map( D => n3032, CK => CLK, Q => n2805, QN =>
                           n2511);
   OUT2_reg_31_inst : DFF_X1 port map( D => n3109, CK => CLK, Q => n2727, QN =>
                           n1315);
   OUT2_reg_30_inst : DFF_X1 port map( D => n3107, CK => CLK, Q => n2729, QN =>
                           n1378);
   OUT2_reg_29_inst : DFF_X1 port map( D => n3105, CK => CLK, Q => n2731, QN =>
                           n1408);
   OUT2_reg_28_inst : DFF_X1 port map( D => n3103, CK => CLK, Q => n2733, QN =>
                           n1438);
   OUT2_reg_27_inst : DFF_X1 port map( D => n3101, CK => CLK, Q => n2735, QN =>
                           n1468);
   OUT2_reg_26_inst : DFF_X1 port map( D => n3099, CK => CLK, Q => n2737, QN =>
                           n1498);
   OUT2_reg_25_inst : DFF_X1 port map( D => n3097, CK => CLK, Q => n2739, QN =>
                           n1528);
   OUT2_reg_24_inst : DFF_X1 port map( D => n3095, CK => CLK, Q => n2741, QN =>
                           n1558);
   OUT1_reg_1_inst : DFF_X1 port map( D => n2986, CK => CLK, Q => n2851, QN => 
                           n4274);
   OUT1_reg_0_inst : DFF_X1 port map( D => n2984, CK => CLK, Q => n2853, QN => 
                           n4295);
   OUT1_reg_23_inst : DFF_X1 port map( D => n3030, CK => CLK, Q => n2807, QN =>
                           n2532);
   OUT1_reg_22_inst : DFF_X1 port map( D => n3028, CK => CLK, Q => n2809, QN =>
                           n2553);
   OUT1_reg_21_inst : DFF_X1 port map( D => n3026, CK => CLK, Q => n2811, QN =>
                           n2574);
   OUT1_reg_20_inst : DFF_X1 port map( D => n3024, CK => CLK, Q => n2813, QN =>
                           n2595);
   OUT1_reg_19_inst : DFF_X1 port map( D => n3022, CK => CLK, Q => n2815, QN =>
                           n2616);
   OUT1_reg_18_inst : DFF_X1 port map( D => n3020, CK => CLK, Q => n2817, QN =>
                           n2637);
   OUT1_reg_17_inst : DFF_X1 port map( D => n3018, CK => CLK, Q => n2819, QN =>
                           n2658);
   OUT1_reg_16_inst : DFF_X1 port map( D => n3016, CK => CLK, Q => n2821, QN =>
                           n2679);
   OUT1_reg_15_inst : DFF_X1 port map( D => n3014, CK => CLK, Q => n2823, QN =>
                           n2700);
   OUT1_reg_14_inst : DFF_X1 port map( D => n3012, CK => CLK, Q => n2825, QN =>
                           n2721);
   OUT1_reg_13_inst : DFF_X1 port map( D => n3010, CK => CLK, Q => n2827, QN =>
                           n2870);
   OUT1_reg_12_inst : DFF_X1 port map( D => n3008, CK => CLK, Q => n2829, QN =>
                           n2891);
   OUT1_reg_11_inst : DFF_X1 port map( D => n3006, CK => CLK, Q => n2831, QN =>
                           n2912);
   OUT1_reg_10_inst : DFF_X1 port map( D => n3004, CK => CLK, Q => n2833, QN =>
                           n2933);
   OUT1_reg_9_inst : DFF_X1 port map( D => n3002, CK => CLK, Q => n2835, QN => 
                           n2954);
   OUT1_reg_8_inst : DFF_X1 port map( D => n3000, CK => CLK, Q => n2837, QN => 
                           n2975);
   OUT1_reg_7_inst : DFF_X1 port map( D => n2998, CK => CLK, Q => n2839, QN => 
                           n4148);
   OUT1_reg_6_inst : DFF_X1 port map( D => n2996, CK => CLK, Q => n2841, QN => 
                           n4169);
   OUT1_reg_5_inst : DFF_X1 port map( D => n2994, CK => CLK, Q => n2843, QN => 
                           n4190);
   OUT1_reg_4_inst : DFF_X1 port map( D => n2992, CK => CLK, Q => n2845, QN => 
                           n4211);
   OUT1_reg_3_inst : DFF_X1 port map( D => n2990, CK => CLK, Q => n2847, QN => 
                           n4232);
   OUT1_reg_2_inst : DFF_X1 port map( D => n2988, CK => CLK, Q => n2849, QN => 
                           n4253);
   OUT2_reg_23_inst : DFF_X1 port map( D => n3093, CK => CLK, Q => n2743, QN =>
                           n1588);
   OUT2_reg_22_inst : DFF_X1 port map( D => n3091, CK => CLK, Q => n2745, QN =>
                           n1618);
   OUT2_reg_19_inst : DFF_X1 port map( D => n3085, CK => CLK, Q => n2751, QN =>
                           n1708);
   OUT2_reg_15_inst : DFF_X1 port map( D => n3077, CK => CLK, Q => n2759, QN =>
                           n1828);
   OUT2_reg_14_inst : DFF_X1 port map( D => n3075, CK => CLK, Q => n2761, QN =>
                           n1858);
   OUT2_reg_11_inst : DFF_X1 port map( D => n3069, CK => CLK, Q => n2767, QN =>
                           n1948);
   OUT2_reg_7_inst : DFF_X1 port map( D => n3061, CK => CLK, Q => n2775, QN => 
                           n2068);
   OUT2_reg_5_inst : DFF_X1 port map( D => n3057, CK => CLK, Q => n2779, QN => 
                           n2128);
   OUT2_reg_3_inst : DFF_X1 port map( D => n3053, CK => CLK, Q => n2783, QN => 
                           n2188);
   OUT2_reg_0_inst : DFF_X1 port map( D => n3047, CK => CLK, Q => n2789, QN => 
                           n2278);
   OUT2_reg_21_inst : DFF_X1 port map( D => n3089, CK => CLK, Q => n2747, QN =>
                           n1648);
   OUT2_reg_20_inst : DFF_X1 port map( D => n3087, CK => CLK, Q => n2749, QN =>
                           n1678);
   OUT2_reg_18_inst : DFF_X1 port map( D => n3083, CK => CLK, Q => n2753, QN =>
                           n1738);
   OUT2_reg_17_inst : DFF_X1 port map( D => n3081, CK => CLK, Q => n2755, QN =>
                           n1768);
   OUT2_reg_16_inst : DFF_X1 port map( D => n3079, CK => CLK, Q => n2757, QN =>
                           n1798);
   OUT2_reg_13_inst : DFF_X1 port map( D => n3073, CK => CLK, Q => n2763, QN =>
                           n1888);
   OUT2_reg_12_inst : DFF_X1 port map( D => n3071, CK => CLK, Q => n2765, QN =>
                           n1918);
   OUT2_reg_10_inst : DFF_X1 port map( D => n3067, CK => CLK, Q => n2769, QN =>
                           n1978);
   OUT2_reg_9_inst : DFF_X1 port map( D => n3065, CK => CLK, Q => n2771, QN => 
                           n2008);
   OUT2_reg_8_inst : DFF_X1 port map( D => n3063, CK => CLK, Q => n2773, QN => 
                           n2038);
   OUT2_reg_6_inst : DFF_X1 port map( D => n3059, CK => CLK, Q => n2777, QN => 
                           n2098);
   OUT2_reg_4_inst : DFF_X1 port map( D => n3055, CK => CLK, Q => n2781, QN => 
                           n2158);
   OUT2_reg_2_inst : DFF_X1 port map( D => n3051, CK => CLK, Q => n2785, QN => 
                           n2218);
   OUT2_reg_1_inst : DFF_X1 port map( D => n3049, CK => CLK, Q => n2787, QN => 
                           n2248);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n4006, CK => CLK, Q => n5267
                           , QN => n128);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n4005, CK => CLK, Q => n5266
                           , QN => n127);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n4004, CK => CLK, Q => n5265
                           , QN => n126);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n4003, CK => CLK, Q => n5264
                           , QN => n125);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n4002, CK => CLK, Q => n5263
                           , QN => n124);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n4001, CK => CLK, Q => n5262
                           , QN => n123);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n4000, CK => CLK, Q => n5261
                           , QN => n122);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n3999, CK => CLK, Q => n5260
                           , QN => n121);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n4038, CK => CLK, Q => n5299
                           , QN => n120);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n4037, CK => CLK, Q => n5298
                           , QN => n119);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n4036, CK => CLK, Q => n5297
                           , QN => n118);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n4035, CK => CLK, Q => n5296
                           , QN => n117);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n4034, CK => CLK, Q => n5295
                           , QN => n116);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n4033, CK => CLK, Q => n5294
                           , QN => n115);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n4032, CK => CLK, Q => n5293
                           , QN => n114);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n4031, CK => CLK, Q => n5292
                           , QN => n113);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n3622, CK => CLK, Q => 
                           n4883, QN => n1351);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n3621, CK => CLK, Q => 
                           n4882, QN => n1395);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n3620, CK => CLK, Q => 
                           n4881, QN => n1425);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n3619, CK => CLK, Q => 
                           n4880, QN => n1455);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n3618, CK => CLK, Q => 
                           n4879, QN => n1485);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n3617, CK => CLK, Q => 
                           n4878, QN => n1515);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n3616, CK => CLK, Q => 
                           n4877, QN => n1545);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n3615, CK => CLK, Q => 
                           n4876, QN => n1575);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n3654, CK => CLK, Q => 
                           n4915, QN => n1353);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n3653, CK => CLK, Q => 
                           n4914, QN => n1396);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n3652, CK => CLK, Q => 
                           n4913, QN => n1426);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n3651, CK => CLK, Q => 
                           n4912, QN => n1456);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n3650, CK => CLK, Q => 
                           n4911, QN => n1486);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n3649, CK => CLK, Q => 
                           n4910, QN => n1516);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n3648, CK => CLK, Q => 
                           n4909, QN => n1546);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n3647, CK => CLK, Q => 
                           n4908, QN => n1576);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n3750, CK => CLK, Q => 
                           n5011, QN => n112);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n3749, CK => CLK, Q => 
                           n5010, QN => n111);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n3748, CK => CLK, Q => 
                           n5009, QN => n110);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n3747, CK => CLK, Q => 
                           n5008, QN => n109);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n3746, CK => CLK, Q => 
                           n5007, QN => n108);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n3745, CK => CLK, Q => 
                           n5006, QN => n107);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n3744, CK => CLK, Q => 
                           n5005, QN => n106);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n3743, CK => CLK, Q => 
                           n5004, QN => n105);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n3878, CK => CLK, Q => n5139
                           , QN => n1360);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n3877, CK => CLK, Q => n5138
                           , QN => n1399);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n3876, CK => CLK, Q => n5137
                           , QN => n1429);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n3875, CK => CLK, Q => n5136
                           , QN => n1459);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n3874, CK => CLK, Q => n5135
                           , QN => n1489);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n3873, CK => CLK, Q => n5134
                           , QN => n1519);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n3872, CK => CLK, Q => n5133
                           , QN => n1549);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n3871, CK => CLK, Q => n5132
                           , QN => n1579);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n3782, CK => CLK, Q => 
                           n5043, QN => n104);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n3781, CK => CLK, Q => 
                           n5042, QN => n103);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n3780, CK => CLK, Q => 
                           n5041, QN => n102);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n3779, CK => CLK, Q => 
                           n5040, QN => n101);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n3778, CK => CLK, Q => 
                           n5039, QN => n100);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n3777, CK => CLK, Q => 
                           n5038, QN => n99);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n3776, CK => CLK, Q => 
                           n5037, QN => n98);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n3775, CK => CLK, Q => 
                           n5036, QN => n97);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n3910, CK => CLK, Q => n5171
                           , QN => n1358);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n3909, CK => CLK, Q => n5170
                           , QN => n1398);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n3908, CK => CLK, Q => n5169
                           , QN => n1428);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n3907, CK => CLK, Q => n5168
                           , QN => n1458);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n3906, CK => CLK, Q => n5167
                           , QN => n1488);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n3905, CK => CLK, Q => n5166
                           , QN => n1518);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n3904, CK => CLK, Q => n5165
                           , QN => n1548);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n3903, CK => CLK, Q => n5164
                           , QN => n1578);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n3998, CK => CLK, Q => n5259
                           , QN => n96);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n3997, CK => CLK, Q => n5258
                           , QN => n95);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n3996, CK => CLK, Q => n5257
                           , QN => n94);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n3995, CK => CLK, Q => n5256
                           , QN => n93);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n3994, CK => CLK, Q => n5255
                           , QN => n92);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n3993, CK => CLK, Q => n5254
                           , QN => n91);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n3992, CK => CLK, Q => n5253
                           , QN => n90);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n3991, CK => CLK, Q => n5252
                           , QN => n89);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n3990, CK => CLK, Q => n5251
                           , QN => n88);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n3989, CK => CLK, Q => n5250
                           , QN => n87);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n3988, CK => CLK, Q => n5249
                           , QN => n86);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n3987, CK => CLK, Q => n5248
                           , QN => n85);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n3986, CK => CLK, Q => n5247
                           , QN => n84);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n3985, CK => CLK, Q => n5246
                           , QN => n83);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n3984, CK => CLK, Q => n5245,
                           QN => n82);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n3983, CK => CLK, Q => n5244,
                           QN => n81);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n3982, CK => CLK, Q => n5243,
                           QN => n80);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n3981, CK => CLK, Q => n5242,
                           QN => n79);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n3980, CK => CLK, Q => n5241,
                           QN => n78);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n3979, CK => CLK, Q => n5240,
                           QN => n77);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n3978, CK => CLK, Q => n5239,
                           QN => n76);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n3977, CK => CLK, Q => n5238,
                           QN => n75);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n3976, CK => CLK, Q => n5237,
                           QN => n74);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n3975, CK => CLK, Q => n5236,
                           QN => n73);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n4030, CK => CLK, Q => n5291
                           , QN => n72);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n4029, CK => CLK, Q => n5290
                           , QN => n71);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n4028, CK => CLK, Q => n5289
                           , QN => n70);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n4027, CK => CLK, Q => n5288
                           , QN => n69);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n4026, CK => CLK, Q => n5287
                           , QN => n68);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n4025, CK => CLK, Q => n5286
                           , QN => n67);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n4024, CK => CLK, Q => n5285
                           , QN => n66);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n4023, CK => CLK, Q => n5284
                           , QN => n65);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n4022, CK => CLK, Q => n5283
                           , QN => n64);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n4021, CK => CLK, Q => n5282
                           , QN => n63);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n4020, CK => CLK, Q => n5281
                           , QN => n62);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n4019, CK => CLK, Q => n5280
                           , QN => n61);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n4018, CK => CLK, Q => n5279
                           , QN => n60);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n4017, CK => CLK, Q => n5278
                           , QN => n59);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n4016, CK => CLK, Q => n5277,
                           QN => n58);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n4015, CK => CLK, Q => n5276,
                           QN => n57);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n4014, CK => CLK, Q => n5275,
                           QN => n56);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n4013, CK => CLK, Q => n5274,
                           QN => n55);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n4012, CK => CLK, Q => n5273,
                           QN => n54);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n4011, CK => CLK, Q => n5272,
                           QN => n53);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n4010, CK => CLK, Q => n5271,
                           QN => n52);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n4009, CK => CLK, Q => n5270,
                           QN => n51);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n4008, CK => CLK, Q => n5269,
                           QN => n50);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n4007, CK => CLK, Q => n5268,
                           QN => n49);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n3614, CK => CLK, Q => 
                           n4875, QN => n1605);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n3613, CK => CLK, Q => 
                           n4874, QN => n1635);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n3612, CK => CLK, Q => 
                           n4873, QN => n1665);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n3611, CK => CLK, Q => 
                           n4872, QN => n1695);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n3610, CK => CLK, Q => 
                           n4871, QN => n1725);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n3609, CK => CLK, Q => 
                           n4870, QN => n1755);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n3608, CK => CLK, Q => 
                           n4869, QN => n1785);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n3607, CK => CLK, Q => 
                           n4868, QN => n1815);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n3606, CK => CLK, Q => 
                           n4867, QN => n1845);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n3605, CK => CLK, Q => 
                           n4866, QN => n1875);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n3604, CK => CLK, Q => 
                           n4865, QN => n1905);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n3603, CK => CLK, Q => 
                           n4864, QN => n1935);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n3602, CK => CLK, Q => 
                           n4863, QN => n1965);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n3601, CK => CLK, Q => 
                           n4862, QN => n1995);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n3600, CK => CLK, Q => n4861
                           , QN => n2025);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n3599, CK => CLK, Q => n4860
                           , QN => n2055);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n3598, CK => CLK, Q => n4859
                           , QN => n2085);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n3597, CK => CLK, Q => n4858
                           , QN => n2115);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n3596, CK => CLK, Q => n4857
                           , QN => n2145);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n3595, CK => CLK, Q => n4856
                           , QN => n2175);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n3594, CK => CLK, Q => n4855
                           , QN => n2205);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n3593, CK => CLK, Q => n4854
                           , QN => n2235);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n3592, CK => CLK, Q => n4853
                           , QN => n2265);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n3591, CK => CLK, Q => n4852
                           , QN => n2307);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n3646, CK => CLK, Q => 
                           n4907, QN => n1606);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n3645, CK => CLK, Q => 
                           n4906, QN => n1636);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n3644, CK => CLK, Q => 
                           n4905, QN => n1666);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n3643, CK => CLK, Q => 
                           n4904, QN => n1696);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n3642, CK => CLK, Q => 
                           n4903, QN => n1726);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n3641, CK => CLK, Q => 
                           n4902, QN => n1756);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n3640, CK => CLK, Q => 
                           n4901, QN => n1786);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n3639, CK => CLK, Q => 
                           n4900, QN => n1816);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n3638, CK => CLK, Q => 
                           n4899, QN => n1846);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n3637, CK => CLK, Q => 
                           n4898, QN => n1876);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n3636, CK => CLK, Q => 
                           n4897, QN => n1906);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n3635, CK => CLK, Q => 
                           n4896, QN => n1936);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n3634, CK => CLK, Q => 
                           n4895, QN => n1966);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n3633, CK => CLK, Q => 
                           n4894, QN => n1996);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n3632, CK => CLK, Q => n4893
                           , QN => n2026);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n3631, CK => CLK, Q => n4892
                           , QN => n2056);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n3630, CK => CLK, Q => n4891
                           , QN => n2086);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n3629, CK => CLK, Q => n4890
                           , QN => n2116);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n3628, CK => CLK, Q => n4889
                           , QN => n2146);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n3627, CK => CLK, Q => n4888
                           , QN => n2176);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n3626, CK => CLK, Q => n4887
                           , QN => n2206);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n3625, CK => CLK, Q => n4886
                           , QN => n2236);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n3624, CK => CLK, Q => n4885
                           , QN => n2266);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n3623, CK => CLK, Q => n4884
                           , QN => n2308);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n3742, CK => CLK, Q => 
                           n5003, QN => n48);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n3741, CK => CLK, Q => 
                           n5002, QN => n47);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n3740, CK => CLK, Q => 
                           n5001, QN => n46);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n3739, CK => CLK, Q => 
                           n5000, QN => n45);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n3738, CK => CLK, Q => 
                           n4999, QN => n44);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n3737, CK => CLK, Q => 
                           n4998, QN => n43);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n3736, CK => CLK, Q => 
                           n4997, QN => n42);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n3735, CK => CLK, Q => 
                           n4996, QN => n41);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n3734, CK => CLK, Q => 
                           n4995, QN => n40);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n3733, CK => CLK, Q => 
                           n4994, QN => n39);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n3732, CK => CLK, Q => 
                           n4993, QN => n38);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n3731, CK => CLK, Q => 
                           n4992, QN => n37);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n3730, CK => CLK, Q => 
                           n4991, QN => n36);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n3729, CK => CLK, Q => 
                           n4990, QN => n35);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n3728, CK => CLK, Q => n4989
                           , QN => n34);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n3727, CK => CLK, Q => n4988
                           , QN => n33);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n3726, CK => CLK, Q => n4987
                           , QN => n32);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n3725, CK => CLK, Q => n4986
                           , QN => n31);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n3724, CK => CLK, Q => n4985
                           , QN => n30);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n3723, CK => CLK, Q => n4984
                           , QN => n29);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n3722, CK => CLK, Q => n4983
                           , QN => n28);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n3721, CK => CLK, Q => n4982
                           , QN => n27);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n3720, CK => CLK, Q => n4981
                           , QN => n26);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n3719, CK => CLK, Q => n4980
                           , QN => n25);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n3870, CK => CLK, Q => n5131
                           , QN => n1609);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n3869, CK => CLK, Q => n5130
                           , QN => n1639);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n3868, CK => CLK, Q => n5129
                           , QN => n1669);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n3867, CK => CLK, Q => n5128
                           , QN => n1699);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n3866, CK => CLK, Q => n5127
                           , QN => n1729);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n3865, CK => CLK, Q => n5126
                           , QN => n1759);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n3864, CK => CLK, Q => n5125
                           , QN => n1789);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n3863, CK => CLK, Q => n5124
                           , QN => n1819);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n3862, CK => CLK, Q => n5123
                           , QN => n1849);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n3861, CK => CLK, Q => n5122
                           , QN => n1879);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n3860, CK => CLK, Q => n5121
                           , QN => n1909);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n3859, CK => CLK, Q => n5120
                           , QN => n1939);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n3858, CK => CLK, Q => n5119
                           , QN => n1969);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n3857, CK => CLK, Q => n5118
                           , QN => n1999);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n3856, CK => CLK, Q => n5117,
                           QN => n2029);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n3855, CK => CLK, Q => n5116,
                           QN => n2059);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n3854, CK => CLK, Q => n5115,
                           QN => n2089);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n3853, CK => CLK, Q => n5114,
                           QN => n2119);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n3852, CK => CLK, Q => n5113,
                           QN => n2149);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n3851, CK => CLK, Q => n5112,
                           QN => n2179);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n3850, CK => CLK, Q => n5111,
                           QN => n2209);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n3849, CK => CLK, Q => n5110,
                           QN => n2239);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n3848, CK => CLK, Q => n5109,
                           QN => n2269);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n3847, CK => CLK, Q => n5108,
                           QN => n2313);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n3774, CK => CLK, Q => 
                           n5035, QN => n24);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n3773, CK => CLK, Q => 
                           n5034, QN => n23);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n3772, CK => CLK, Q => 
                           n5033, QN => n22);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n3771, CK => CLK, Q => 
                           n5032, QN => n21);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n3770, CK => CLK, Q => 
                           n5031, QN => n20);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n3769, CK => CLK, Q => 
                           n5030, QN => n19);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n3768, CK => CLK, Q => 
                           n5029, QN => n18);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n3767, CK => CLK, Q => 
                           n5028, QN => n17);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n3766, CK => CLK, Q => 
                           n5027, QN => n16);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n3765, CK => CLK, Q => 
                           n5026, QN => n15);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n3764, CK => CLK, Q => 
                           n5025, QN => n14);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n3763, CK => CLK, Q => 
                           n5024, QN => n13);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n3762, CK => CLK, Q => 
                           n5023, QN => n12);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n3761, CK => CLK, Q => 
                           n5022, QN => n11);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n3760, CK => CLK, Q => n5021
                           , QN => n10);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n3759, CK => CLK, Q => n5020
                           , QN => n9);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n3758, CK => CLK, Q => n5019
                           , QN => n8);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n3757, CK => CLK, Q => n5018
                           , QN => n7);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n3756, CK => CLK, Q => n5017
                           , QN => n6);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n3755, CK => CLK, Q => n5016
                           , QN => n5);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n3754, CK => CLK, Q => n5015
                           , QN => n4);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n3753, CK => CLK, Q => n5014
                           , QN => n3);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n3752, CK => CLK, Q => n5013
                           , QN => n2);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n3751, CK => CLK, Q => n5012
                           , QN => n1);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n3902, CK => CLK, Q => n5163
                           , QN => n1608);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n3901, CK => CLK, Q => n5162
                           , QN => n1638);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n3900, CK => CLK, Q => n5161
                           , QN => n1668);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n3899, CK => CLK, Q => n5160
                           , QN => n1698);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n3898, CK => CLK, Q => n5159
                           , QN => n1728);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n3897, CK => CLK, Q => n5158
                           , QN => n1758);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n3896, CK => CLK, Q => n5157
                           , QN => n1788);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n3895, CK => CLK, Q => n5156
                           , QN => n1818);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n3894, CK => CLK, Q => n5155
                           , QN => n1848);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n3893, CK => CLK, Q => n5154
                           , QN => n1878);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n3892, CK => CLK, Q => n5153
                           , QN => n1908);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n3891, CK => CLK, Q => n5152
                           , QN => n1938);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n3890, CK => CLK, Q => n5151
                           , QN => n1968);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n3889, CK => CLK, Q => n5150
                           , QN => n1998);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n3888, CK => CLK, Q => n5149,
                           QN => n2028);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n3887, CK => CLK, Q => n5148,
                           QN => n2058);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n3886, CK => CLK, Q => n5147,
                           QN => n2088);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n3885, CK => CLK, Q => n5146,
                           QN => n2118);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n3884, CK => CLK, Q => n5145,
                           QN => n2148);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n3883, CK => CLK, Q => n5144,
                           QN => n2178);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n3882, CK => CLK, Q => n5143,
                           QN => n2208);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n3881, CK => CLK, Q => n5142,
                           QN => n2238);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n3880, CK => CLK, Q => n5141,
                           QN => n2268);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n3879, CK => CLK, Q => n5140,
                           QN => n2312);
   U3 : BUF_X1 port map( A => n2334, Z => n610);
   U4 : BUF_X1 port map( A => n2334, Z => n611);
   U5 : BUF_X1 port map( A => n1319, Z => n508);
   U6 : BUF_X1 port map( A => n1319, Z => n509);
   U7 : BUF_X1 port map( A => n441, Z => n442);
   U8 : BUF_X1 port map( A => n441, Z => n443);
   U9 : BUF_X1 port map( A => n284, Z => n285);
   U10 : BUF_X1 port map( A => n284, Z => n286);
   U11 : BUF_X1 port map( A => n441, Z => n444);
   U12 : BUF_X1 port map( A => n284, Z => n287);
   U13 : BUF_X1 port map( A => n2334, Z => n612);
   U14 : BUF_X1 port map( A => n1319, Z => n510);
   U15 : BUF_X1 port map( A => n2349, Z => n637);
   U16 : BUF_X1 port map( A => n2349, Z => n638);
   U17 : BUF_X1 port map( A => n1334, Z => n535);
   U18 : BUF_X1 port map( A => n1334, Z => n536);
   U19 : BUF_X1 port map( A => n2349, Z => n639);
   U20 : BUF_X1 port map( A => n1334, Z => n537);
   U21 : BUF_X1 port map( A => n257, Z => n261);
   U22 : BUF_X1 port map( A => n257, Z => n260);
   U23 : BUF_X1 port map( A => n257, Z => n262);
   U24 : BUF_X1 port map( A => n257, Z => n263);
   U25 : BUF_X1 port map( A => n257, Z => n264);
   U26 : BUF_X1 port map( A => n257, Z => n265);
   U27 : BUF_X1 port map( A => n258, Z => n269);
   U28 : BUF_X1 port map( A => n258, Z => n266);
   U29 : BUF_X1 port map( A => n258, Z => n267);
   U30 : BUF_X1 port map( A => n258, Z => n268);
   U31 : BUF_X1 port map( A => n258, Z => n270);
   U32 : BUF_X1 port map( A => n258, Z => n271);
   U33 : BUF_X1 port map( A => n259, Z => n273);
   U34 : BUF_X1 port map( A => n259, Z => n274);
   U35 : BUF_X1 port map( A => n259, Z => n272);
   U36 : BUF_X1 port map( A => n259, Z => n275);
   U37 : BUF_X1 port map( A => n501, Z => n502);
   U38 : BUF_X1 port map( A => n501, Z => n503);
   U39 : BUF_X1 port map( A => n497, Z => n498);
   U40 : BUF_X1 port map( A => n497, Z => n499);
   U41 : BUF_X1 port map( A => n493, Z => n494);
   U42 : BUF_X1 port map( A => n493, Z => n495);
   U43 : BUF_X1 port map( A => n489, Z => n490);
   U44 : BUF_X1 port map( A => n489, Z => n491);
   U45 : BUF_X1 port map( A => n485, Z => n486);
   U46 : BUF_X1 port map( A => n485, Z => n487);
   U47 : BUF_X1 port map( A => n481, Z => n482);
   U48 : BUF_X1 port map( A => n481, Z => n483);
   U49 : BUF_X1 port map( A => n477, Z => n478);
   U50 : BUF_X1 port map( A => n477, Z => n479);
   U51 : BUF_X1 port map( A => n473, Z => n474);
   U52 : BUF_X1 port map( A => n473, Z => n475);
   U53 : BUF_X1 port map( A => n469, Z => n470);
   U54 : BUF_X1 port map( A => n469, Z => n471);
   U55 : BUF_X1 port map( A => n465, Z => n466);
   U56 : BUF_X1 port map( A => n465, Z => n467);
   U57 : BUF_X1 port map( A => n461, Z => n462);
   U58 : BUF_X1 port map( A => n461, Z => n463);
   U59 : BUF_X1 port map( A => n457, Z => n458);
   U60 : BUF_X1 port map( A => n457, Z => n459);
   U61 : BUF_X1 port map( A => n453, Z => n454);
   U62 : BUF_X1 port map( A => n453, Z => n455);
   U63 : BUF_X1 port map( A => n449, Z => n450);
   U64 : BUF_X1 port map( A => n449, Z => n451);
   U65 : BUF_X1 port map( A => n445, Z => n446);
   U66 : BUF_X1 port map( A => n445, Z => n447);
   U67 : BUF_X1 port map( A => n437, Z => n438);
   U68 : BUF_X1 port map( A => n437, Z => n439);
   U69 : BUF_X1 port map( A => n433, Z => n434);
   U70 : BUF_X1 port map( A => n433, Z => n435);
   U71 : BUF_X1 port map( A => n429, Z => n430);
   U72 : BUF_X1 port map( A => n429, Z => n431);
   U73 : BUF_X1 port map( A => n425, Z => n426);
   U74 : BUF_X1 port map( A => n425, Z => n427);
   U75 : BUF_X1 port map( A => n421, Z => n422);
   U76 : BUF_X1 port map( A => n421, Z => n423);
   U77 : BUF_X1 port map( A => n417, Z => n418);
   U78 : BUF_X1 port map( A => n417, Z => n419);
   U79 : BUF_X1 port map( A => n413, Z => n414);
   U80 : BUF_X1 port map( A => n413, Z => n415);
   U81 : BUF_X1 port map( A => n409, Z => n410);
   U82 : BUF_X1 port map( A => n409, Z => n411);
   U83 : BUF_X1 port map( A => n405, Z => n406);
   U84 : BUF_X1 port map( A => n405, Z => n407);
   U85 : BUF_X1 port map( A => n401, Z => n402);
   U86 : BUF_X1 port map( A => n401, Z => n403);
   U87 : BUF_X1 port map( A => n397, Z => n398);
   U88 : BUF_X1 port map( A => n397, Z => n399);
   U89 : BUF_X1 port map( A => n393, Z => n394);
   U90 : BUF_X1 port map( A => n393, Z => n395);
   U91 : BUF_X1 port map( A => n389, Z => n390);
   U92 : BUF_X1 port map( A => n389, Z => n391);
   U93 : BUF_X1 port map( A => n385, Z => n386);
   U94 : BUF_X1 port map( A => n385, Z => n387);
   U95 : BUF_X1 port map( A => n381, Z => n382);
   U96 : BUF_X1 port map( A => n381, Z => n383);
   U97 : BUF_X1 port map( A => n501, Z => n504);
   U98 : BUF_X1 port map( A => n497, Z => n500);
   U99 : BUF_X1 port map( A => n493, Z => n496);
   U100 : BUF_X1 port map( A => n489, Z => n492);
   U101 : BUF_X1 port map( A => n485, Z => n488);
   U102 : BUF_X1 port map( A => n481, Z => n484);
   U103 : BUF_X1 port map( A => n477, Z => n480);
   U104 : BUF_X1 port map( A => n473, Z => n476);
   U105 : BUF_X1 port map( A => n469, Z => n472);
   U106 : BUF_X1 port map( A => n465, Z => n468);
   U107 : BUF_X1 port map( A => n461, Z => n464);
   U108 : BUF_X1 port map( A => n457, Z => n460);
   U109 : BUF_X1 port map( A => n453, Z => n456);
   U110 : BUF_X1 port map( A => n449, Z => n452);
   U111 : BUF_X1 port map( A => n445, Z => n448);
   U112 : BUF_X1 port map( A => n437, Z => n440);
   U113 : BUF_X1 port map( A => n433, Z => n436);
   U114 : BUF_X1 port map( A => n429, Z => n432);
   U115 : BUF_X1 port map( A => n425, Z => n428);
   U116 : BUF_X1 port map( A => n421, Z => n424);
   U117 : BUF_X1 port map( A => n417, Z => n420);
   U118 : BUF_X1 port map( A => n413, Z => n416);
   U119 : BUF_X1 port map( A => n409, Z => n412);
   U120 : BUF_X1 port map( A => n405, Z => n408);
   U121 : BUF_X1 port map( A => n401, Z => n404);
   U122 : BUF_X1 port map( A => n397, Z => n400);
   U123 : BUF_X1 port map( A => n393, Z => n396);
   U124 : BUF_X1 port map( A => n389, Z => n392);
   U125 : BUF_X1 port map( A => n385, Z => n388);
   U126 : BUF_X1 port map( A => n381, Z => n384);
   U127 : BUF_X1 port map( A => n709, Z => n710);
   U128 : BUF_X1 port map( A => n709, Z => n711);
   U129 : BUF_X1 port map( A => n277, Z => n278);
   U130 : BUF_X1 port map( A => n277, Z => n279);
   U131 : BUF_X1 port map( A => n709, Z => n712);
   U132 : BUF_X1 port map( A => n277, Z => n280);
   U133 : BUF_X1 port map( A => n813, Z => n379);
   U134 : BUF_X1 port map( A => n811, Z => n376);
   U135 : BUF_X1 port map( A => n809, Z => n373);
   U136 : BUF_X1 port map( A => n807, Z => n370);
   U137 : BUF_X1 port map( A => n805, Z => n367);
   U138 : BUF_X1 port map( A => n803, Z => n364);
   U139 : BUF_X1 port map( A => n801, Z => n361);
   U140 : BUF_X1 port map( A => n799, Z => n358);
   U141 : BUF_X1 port map( A => n797, Z => n355);
   U142 : BUF_X1 port map( A => n795, Z => n352);
   U143 : BUF_X1 port map( A => n793, Z => n349);
   U144 : BUF_X1 port map( A => n791, Z => n346);
   U145 : BUF_X1 port map( A => n789, Z => n343);
   U146 : BUF_X1 port map( A => n787, Z => n340);
   U147 : BUF_X1 port map( A => n785, Z => n337);
   U148 : BUF_X1 port map( A => n783, Z => n334);
   U149 : BUF_X1 port map( A => n781, Z => n331);
   U150 : BUF_X1 port map( A => n779, Z => n328);
   U151 : BUF_X1 port map( A => n777, Z => n325);
   U152 : BUF_X1 port map( A => n775, Z => n322);
   U153 : BUF_X1 port map( A => n773, Z => n319);
   U154 : BUF_X1 port map( A => n771, Z => n316);
   U155 : BUF_X1 port map( A => n769, Z => n313);
   U156 : BUF_X1 port map( A => n767, Z => n310);
   U157 : BUF_X1 port map( A => n765, Z => n307);
   U158 : BUF_X1 port map( A => n763, Z => n304);
   U159 : BUF_X1 port map( A => n761, Z => n301);
   U160 : BUF_X1 port map( A => n759, Z => n298);
   U161 : BUF_X1 port map( A => n757, Z => n295);
   U162 : BUF_X1 port map( A => n755, Z => n292);
   U163 : BUF_X1 port map( A => n753, Z => n289);
   U164 : BUF_X1 port map( A => n750, Z => n282);
   U165 : BUF_X1 port map( A => n813, Z => n378);
   U166 : BUF_X1 port map( A => n811, Z => n375);
   U167 : BUF_X1 port map( A => n809, Z => n372);
   U168 : BUF_X1 port map( A => n807, Z => n369);
   U169 : BUF_X1 port map( A => n805, Z => n366);
   U170 : BUF_X1 port map( A => n803, Z => n363);
   U171 : BUF_X1 port map( A => n801, Z => n360);
   U172 : BUF_X1 port map( A => n799, Z => n357);
   U173 : BUF_X1 port map( A => n797, Z => n354);
   U174 : BUF_X1 port map( A => n795, Z => n351);
   U175 : BUF_X1 port map( A => n793, Z => n348);
   U176 : BUF_X1 port map( A => n791, Z => n345);
   U177 : BUF_X1 port map( A => n789, Z => n342);
   U178 : BUF_X1 port map( A => n787, Z => n339);
   U179 : BUF_X1 port map( A => n785, Z => n336);
   U180 : BUF_X1 port map( A => n783, Z => n333);
   U181 : BUF_X1 port map( A => n781, Z => n330);
   U182 : BUF_X1 port map( A => n779, Z => n327);
   U183 : BUF_X1 port map( A => n777, Z => n324);
   U184 : BUF_X1 port map( A => n775, Z => n321);
   U185 : BUF_X1 port map( A => n773, Z => n318);
   U186 : BUF_X1 port map( A => n771, Z => n315);
   U187 : BUF_X1 port map( A => n769, Z => n312);
   U188 : BUF_X1 port map( A => n767, Z => n309);
   U189 : BUF_X1 port map( A => n765, Z => n306);
   U190 : BUF_X1 port map( A => n763, Z => n303);
   U191 : BUF_X1 port map( A => n761, Z => n300);
   U192 : BUF_X1 port map( A => n759, Z => n297);
   U193 : BUF_X1 port map( A => n757, Z => n294);
   U194 : BUF_X1 port map( A => n755, Z => n291);
   U195 : BUF_X1 port map( A => n753, Z => n288);
   U196 : BUF_X1 port map( A => n750, Z => n281);
   U197 : BUF_X1 port map( A => n813, Z => n380);
   U198 : BUF_X1 port map( A => n811, Z => n377);
   U199 : BUF_X1 port map( A => n809, Z => n374);
   U200 : BUF_X1 port map( A => n807, Z => n371);
   U201 : BUF_X1 port map( A => n805, Z => n368);
   U202 : BUF_X1 port map( A => n803, Z => n365);
   U203 : BUF_X1 port map( A => n801, Z => n362);
   U204 : BUF_X1 port map( A => n799, Z => n359);
   U205 : BUF_X1 port map( A => n797, Z => n356);
   U206 : BUF_X1 port map( A => n795, Z => n353);
   U207 : BUF_X1 port map( A => n793, Z => n350);
   U208 : BUF_X1 port map( A => n791, Z => n347);
   U209 : BUF_X1 port map( A => n789, Z => n344);
   U210 : BUF_X1 port map( A => n787, Z => n341);
   U211 : BUF_X1 port map( A => n785, Z => n338);
   U212 : BUF_X1 port map( A => n783, Z => n335);
   U213 : BUF_X1 port map( A => n781, Z => n332);
   U214 : BUF_X1 port map( A => n779, Z => n329);
   U215 : BUF_X1 port map( A => n777, Z => n326);
   U216 : BUF_X1 port map( A => n775, Z => n323);
   U217 : BUF_X1 port map( A => n773, Z => n320);
   U218 : BUF_X1 port map( A => n771, Z => n317);
   U219 : BUF_X1 port map( A => n769, Z => n314);
   U220 : BUF_X1 port map( A => n767, Z => n311);
   U221 : BUF_X1 port map( A => n765, Z => n308);
   U222 : BUF_X1 port map( A => n763, Z => n305);
   U223 : BUF_X1 port map( A => n761, Z => n302);
   U224 : BUF_X1 port map( A => n759, Z => n299);
   U225 : BUF_X1 port map( A => n757, Z => n296);
   U226 : BUF_X1 port map( A => n755, Z => n293);
   U227 : BUF_X1 port map( A => n753, Z => n290);
   U228 : BUF_X1 port map( A => n750, Z => n283);
   U229 : BUF_X1 port map( A => n1066, Z => n441);
   U230 : BUF_X1 port map( A => n751, Z => n284);
   U231 : BUF_X1 port map( A => n2345, Z => n628);
   U232 : BUF_X1 port map( A => n2340, Z => n616);
   U233 : BUF_X1 port map( A => n2345, Z => n629);
   U234 : BUF_X1 port map( A => n2340, Z => n617);
   U235 : BUF_X1 port map( A => n1330, Z => n526);
   U236 : BUF_X1 port map( A => n1325, Z => n514);
   U237 : BUF_X1 port map( A => n1330, Z => n527);
   U238 : BUF_X1 port map( A => n1325, Z => n515);
   U239 : BUF_X1 port map( A => n2374, Z => n688);
   U240 : BUF_X1 port map( A => n2369, Z => n676);
   U241 : BUF_X1 port map( A => n2364, Z => n664);
   U242 : BUF_X1 port map( A => n2379, Z => n700);
   U243 : BUF_X1 port map( A => n2350, Z => n640);
   U244 : BUF_X1 port map( A => n2355, Z => n652);
   U245 : BUF_X1 port map( A => n2374, Z => n689);
   U246 : BUF_X1 port map( A => n2369, Z => n677);
   U247 : BUF_X1 port map( A => n2364, Z => n665);
   U248 : BUF_X1 port map( A => n2379, Z => n701);
   U249 : BUF_X1 port map( A => n2350, Z => n641);
   U250 : BUF_X1 port map( A => n2355, Z => n653);
   U251 : BUF_X1 port map( A => n1363, Z => n586);
   U252 : BUF_X1 port map( A => n1356, Z => n574);
   U253 : BUF_X1 port map( A => n1349, Z => n562);
   U254 : BUF_X1 port map( A => n1370, Z => n598);
   U255 : BUF_X1 port map( A => n1335, Z => n538);
   U256 : BUF_X1 port map( A => n1340, Z => n550);
   U257 : BUF_X1 port map( A => n1363, Z => n587);
   U258 : BUF_X1 port map( A => n1356, Z => n575);
   U259 : BUF_X1 port map( A => n1349, Z => n563);
   U260 : BUF_X1 port map( A => n1370, Z => n599);
   U261 : BUF_X1 port map( A => n1335, Z => n539);
   U262 : BUF_X1 port map( A => n1340, Z => n551);
   U263 : BUF_X1 port map( A => n2372, Z => n682);
   U264 : BUF_X1 port map( A => n2382, Z => n706);
   U265 : BUF_X1 port map( A => n2353, Z => n646);
   U266 : BUF_X1 port map( A => n2372, Z => n683);
   U267 : BUF_X1 port map( A => n2382, Z => n707);
   U268 : BUF_X1 port map( A => n2353, Z => n647);
   U269 : BUF_X1 port map( A => n1361, Z => n580);
   U270 : BUF_X1 port map( A => n1375, Z => n604);
   U271 : BUF_X1 port map( A => n1338, Z => n544);
   U272 : BUF_X1 port map( A => n1361, Z => n581);
   U273 : BUF_X1 port map( A => n1375, Z => n605);
   U274 : BUF_X1 port map( A => n1338, Z => n545);
   U275 : BUF_X1 port map( A => n2358, Z => n658);
   U276 : BUF_X1 port map( A => n2358, Z => n659);
   U277 : BUF_X1 port map( A => n1343, Z => n556);
   U278 : BUF_X1 port map( A => n1343, Z => n557);
   U279 : BUF_X1 port map( A => n2377, Z => n694);
   U280 : BUF_X1 port map( A => n2367, Z => n670);
   U281 : BUF_X1 port map( A => n2348, Z => n634);
   U282 : BUF_X1 port map( A => n2343, Z => n622);
   U283 : BUF_X1 port map( A => n2377, Z => n695);
   U284 : BUF_X1 port map( A => n2367, Z => n671);
   U285 : BUF_X1 port map( A => n2348, Z => n635);
   U286 : BUF_X1 port map( A => n2343, Z => n623);
   U287 : BUF_X1 port map( A => n1368, Z => n592);
   U288 : BUF_X1 port map( A => n1354, Z => n568);
   U289 : BUF_X1 port map( A => n1333, Z => n532);
   U290 : BUF_X1 port map( A => n1328, Z => n520);
   U291 : BUF_X1 port map( A => n1368, Z => n593);
   U292 : BUF_X1 port map( A => n1354, Z => n569);
   U293 : BUF_X1 port map( A => n1333, Z => n533);
   U294 : BUF_X1 port map( A => n1328, Z => n521);
   U295 : BUF_X1 port map( A => n2371, Z => n679);
   U296 : BUF_X1 port map( A => n2381, Z => n703);
   U297 : BUF_X1 port map( A => n2352, Z => n643);
   U298 : BUF_X1 port map( A => n2371, Z => n680);
   U299 : BUF_X1 port map( A => n2381, Z => n704);
   U300 : BUF_X1 port map( A => n2352, Z => n644);
   U301 : BUF_X1 port map( A => n1359, Z => n577);
   U302 : BUF_X1 port map( A => n1373, Z => n601);
   U303 : BUF_X1 port map( A => n1337, Z => n541);
   U304 : BUF_X1 port map( A => n1359, Z => n578);
   U305 : BUF_X1 port map( A => n1373, Z => n602);
   U306 : BUF_X1 port map( A => n1337, Z => n542);
   U307 : BUF_X1 port map( A => n2357, Z => n655);
   U308 : BUF_X1 port map( A => n2357, Z => n656);
   U309 : BUF_X1 port map( A => n1342, Z => n553);
   U310 : BUF_X1 port map( A => n1342, Z => n554);
   U311 : BUF_X1 port map( A => n2376, Z => n691);
   U312 : BUF_X1 port map( A => n2366, Z => n667);
   U313 : BUF_X1 port map( A => n2342, Z => n619);
   U314 : BUF_X1 port map( A => n2376, Z => n692);
   U315 : BUF_X1 port map( A => n2366, Z => n668);
   U316 : BUF_X1 port map( A => n2342, Z => n620);
   U317 : BUF_X1 port map( A => n1366, Z => n589);
   U318 : BUF_X1 port map( A => n1352, Z => n565);
   U319 : BUF_X1 port map( A => n1327, Z => n517);
   U320 : BUF_X1 port map( A => n1366, Z => n590);
   U321 : BUF_X1 port map( A => n1352, Z => n566);
   U322 : BUF_X1 port map( A => n1327, Z => n518);
   U323 : BUF_X1 port map( A => n2347, Z => n631);
   U324 : BUF_X1 port map( A => n2347, Z => n632);
   U325 : BUF_X1 port map( A => n1332, Z => n529);
   U326 : BUF_X1 port map( A => n1332, Z => n530);
   U327 : BUF_X1 port map( A => n2373, Z => n685);
   U328 : BUF_X1 port map( A => n2363, Z => n661);
   U329 : BUF_X1 port map( A => n2344, Z => n625);
   U330 : BUF_X1 port map( A => n2339, Z => n613);
   U331 : BUF_X1 port map( A => n2373, Z => n686);
   U332 : BUF_X1 port map( A => n2363, Z => n662);
   U333 : BUF_X1 port map( A => n2344, Z => n626);
   U334 : BUF_X1 port map( A => n2339, Z => n614);
   U335 : BUF_X1 port map( A => n1362, Z => n583);
   U336 : BUF_X1 port map( A => n1348, Z => n559);
   U337 : BUF_X1 port map( A => n1329, Z => n523);
   U338 : BUF_X1 port map( A => n1324, Z => n511);
   U339 : BUF_X1 port map( A => n1362, Z => n584);
   U340 : BUF_X1 port map( A => n1348, Z => n560);
   U341 : BUF_X1 port map( A => n1329, Z => n524);
   U342 : BUF_X1 port map( A => n1324, Z => n512);
   U343 : BUF_X1 port map( A => n2368, Z => n673);
   U344 : BUF_X1 port map( A => n2378, Z => n697);
   U345 : BUF_X1 port map( A => n2354, Z => n649);
   U346 : BUF_X1 port map( A => n2368, Z => n674);
   U347 : BUF_X1 port map( A => n2378, Z => n698);
   U348 : BUF_X1 port map( A => n2354, Z => n650);
   U349 : BUF_X1 port map( A => n1355, Z => n571);
   U350 : BUF_X1 port map( A => n1369, Z => n595);
   U351 : BUF_X1 port map( A => n1339, Z => n547);
   U352 : BUF_X1 port map( A => n1355, Z => n572);
   U353 : BUF_X1 port map( A => n1369, Z => n596);
   U354 : BUF_X1 port map( A => n1339, Z => n548);
   U355 : BUF_X1 port map( A => n2345, Z => n630);
   U356 : BUF_X1 port map( A => n2340, Z => n618);
   U357 : BUF_X1 port map( A => n1330, Z => n528);
   U358 : BUF_X1 port map( A => n1325, Z => n516);
   U359 : BUF_X1 port map( A => n2374, Z => n690);
   U360 : BUF_X1 port map( A => n2369, Z => n678);
   U361 : BUF_X1 port map( A => n2364, Z => n666);
   U362 : BUF_X1 port map( A => n2379, Z => n702);
   U363 : BUF_X1 port map( A => n2350, Z => n642);
   U364 : BUF_X1 port map( A => n1356, Z => n576);
   U365 : BUF_X1 port map( A => n1349, Z => n564);
   U366 : BUF_X1 port map( A => n2355, Z => n654);
   U367 : BUF_X1 port map( A => n1363, Z => n588);
   U368 : BUF_X1 port map( A => n1370, Z => n600);
   U369 : BUF_X1 port map( A => n1335, Z => n540);
   U370 : BUF_X1 port map( A => n1340, Z => n552);
   U371 : BUF_X1 port map( A => n2372, Z => n684);
   U372 : BUF_X1 port map( A => n2382, Z => n708);
   U373 : BUF_X1 port map( A => n2353, Z => n648);
   U374 : BUF_X1 port map( A => n1361, Z => n582);
   U375 : BUF_X1 port map( A => n1375, Z => n606);
   U376 : BUF_X1 port map( A => n1338, Z => n546);
   U377 : BUF_X1 port map( A => n2358, Z => n660);
   U378 : BUF_X1 port map( A => n1343, Z => n558);
   U379 : BUF_X1 port map( A => n2377, Z => n696);
   U380 : BUF_X1 port map( A => n2367, Z => n672);
   U381 : BUF_X1 port map( A => n2343, Z => n624);
   U382 : BUF_X1 port map( A => n1368, Z => n594);
   U383 : BUF_X1 port map( A => n1354, Z => n570);
   U384 : BUF_X1 port map( A => n1328, Z => n522);
   U385 : BUF_X1 port map( A => n2348, Z => n636);
   U386 : BUF_X1 port map( A => n1333, Z => n534);
   U387 : BUF_X1 port map( A => n2371, Z => n681);
   U388 : BUF_X1 port map( A => n2381, Z => n705);
   U389 : BUF_X1 port map( A => n2352, Z => n645);
   U390 : BUF_X1 port map( A => n1359, Z => n579);
   U391 : BUF_X1 port map( A => n1373, Z => n603);
   U392 : BUF_X1 port map( A => n1337, Z => n543);
   U393 : BUF_X1 port map( A => n2357, Z => n657);
   U394 : BUF_X1 port map( A => n1342, Z => n555);
   U395 : BUF_X1 port map( A => n2376, Z => n693);
   U396 : BUF_X1 port map( A => n2366, Z => n669);
   U397 : BUF_X1 port map( A => n2342, Z => n621);
   U398 : BUF_X1 port map( A => n1366, Z => n591);
   U399 : BUF_X1 port map( A => n1352, Z => n567);
   U400 : BUF_X1 port map( A => n1327, Z => n519);
   U401 : BUF_X1 port map( A => n2347, Z => n633);
   U402 : BUF_X1 port map( A => n1332, Z => n531);
   U403 : BUF_X1 port map( A => n2363, Z => n663);
   U404 : BUF_X1 port map( A => n1348, Z => n561);
   U405 : BUF_X1 port map( A => n2373, Z => n687);
   U406 : BUF_X1 port map( A => n2344, Z => n627);
   U407 : BUF_X1 port map( A => n2339, Z => n615);
   U408 : BUF_X1 port map( A => n1362, Z => n585);
   U409 : BUF_X1 port map( A => n1329, Z => n525);
   U410 : BUF_X1 port map( A => n1324, Z => n513);
   U411 : BUF_X1 port map( A => n2368, Z => n675);
   U412 : BUF_X1 port map( A => n2378, Z => n699);
   U413 : BUF_X1 port map( A => n2354, Z => n651);
   U414 : BUF_X1 port map( A => n1355, Z => n573);
   U415 : BUF_X1 port map( A => n1369, Z => n597);
   U416 : BUF_X1 port map( A => n1339, Z => n549);
   U417 : BUF_X1 port map( A => n2329, Z => n608);
   U418 : BUF_X1 port map( A => n2329, Z => n607);
   U419 : BUF_X1 port map( A => n1314, Z => n506);
   U420 : BUF_X1 port map( A => n1314, Z => n505);
   U421 : BUF_X1 port map( A => n2329, Z => n609);
   U422 : BUF_X1 port map( A => n1314, Z => n507);
   U423 : BUF_X1 port map( A => n713, Z => n257);
   U424 : BUF_X1 port map( A => n713, Z => n258);
   U425 : BUF_X1 port map( A => n713, Z => n259);
   U426 : BUF_X1 port map( A => n1312, Z => n501);
   U427 : BUF_X1 port map( A => n1279, Z => n497);
   U428 : BUF_X1 port map( A => n1277, Z => n493);
   U429 : BUF_X1 port map( A => n1273, Z => n489);
   U430 : BUF_X1 port map( A => n1241, Z => n485);
   U431 : BUF_X1 port map( A => n1208, Z => n481);
   U432 : BUF_X1 port map( A => n1206, Z => n477);
   U433 : BUF_X1 port map( A => n1204, Z => n473);
   U434 : BUF_X1 port map( A => n1203, Z => n469);
   U435 : BUF_X1 port map( A => n1202, Z => n465);
   U436 : BUF_X1 port map( A => n1170, Z => n461);
   U437 : BUF_X1 port map( A => n1136, Z => n457);
   U438 : BUF_X1 port map( A => n1133, Z => n453);
   U439 : BUF_X1 port map( A => n1132, Z => n449);
   U440 : BUF_X1 port map( A => n1100, Z => n445);
   U441 : BUF_X1 port map( A => n1063, Z => n437);
   U442 : BUF_X1 port map( A => n1062, Z => n433);
   U443 : BUF_X1 port map( A => n1030, Z => n429);
   U444 : BUF_X1 port map( A => n996, Z => n425);
   U445 : BUF_X1 port map( A => n994, Z => n421);
   U446 : BUF_X1 port map( A => n993, Z => n417);
   U447 : BUF_X1 port map( A => n961, Z => n413);
   U448 : BUF_X1 port map( A => n927, Z => n409);
   U449 : BUF_X1 port map( A => n925, Z => n405);
   U450 : BUF_X1 port map( A => n924, Z => n401);
   U451 : BUF_X1 port map( A => n892, Z => n397);
   U452 : BUF_X1 port map( A => n858, Z => n393);
   U453 : BUF_X1 port map( A => n852, Z => n389);
   U454 : BUF_X1 port map( A => n850, Z => n385);
   U455 : BUF_X1 port map( A => n817, Z => n381);
   U456 : BUF_X1 port map( A => n2384, Z => n709);
   U457 : BUF_X1 port map( A => n715, Z => n277);
   U458 : CLKBUF_X1 port map( A => n259, Z => n276);
   U459 : OAI21_X1 port map( B1 => n268, B2 => n714, A => n280, ZN => n4134);
   U460 : OAI21_X1 port map( B1 => n265, B2 => n716, A => n280, ZN => n4133);
   U461 : OAI21_X1 port map( B1 => n265, B2 => n717, A => n280, ZN => n4132);
   U462 : OAI21_X1 port map( B1 => n267, B2 => n718, A => n280, ZN => n4131);
   U463 : OAI21_X1 port map( B1 => n267, B2 => n719, A => n280, ZN => n4130);
   U464 : OAI21_X1 port map( B1 => n265, B2 => n720, A => n280, ZN => n4129);
   U465 : OAI21_X1 port map( B1 => n265, B2 => n721, A => n280, ZN => n4128);
   U466 : OAI21_X1 port map( B1 => n265, B2 => n722, A => n280, ZN => n4127);
   U467 : OAI21_X1 port map( B1 => n267, B2 => n723, A => n279, ZN => n4126);
   U468 : OAI21_X1 port map( B1 => n265, B2 => n724, A => n279, ZN => n4125);
   U469 : OAI21_X1 port map( B1 => n267, B2 => n725, A => n279, ZN => n4124);
   U470 : OAI21_X1 port map( B1 => n268, B2 => n726, A => n279, ZN => n4123);
   U471 : OAI21_X1 port map( B1 => n266, B2 => n727, A => n279, ZN => n4122);
   U472 : OAI21_X1 port map( B1 => n266, B2 => n728, A => n279, ZN => n4121);
   U473 : OAI21_X1 port map( B1 => n266, B2 => n729, A => n279, ZN => n4120);
   U474 : OAI21_X1 port map( B1 => n266, B2 => n730, A => n279, ZN => n4119);
   U475 : OAI21_X1 port map( B1 => n267, B2 => n731, A => n279, ZN => n4118);
   U476 : OAI21_X1 port map( B1 => n266, B2 => n732, A => n279, ZN => n4117);
   U477 : OAI21_X1 port map( B1 => n266, B2 => n733, A => n279, ZN => n4116);
   U478 : OAI21_X1 port map( B1 => n267, B2 => n734, A => n279, ZN => n4115);
   U479 : OAI21_X1 port map( B1 => n266, B2 => n735, A => n278, ZN => n4114);
   U480 : OAI21_X1 port map( B1 => n266, B2 => n736, A => n278, ZN => n4113);
   U481 : OAI21_X1 port map( B1 => n267, B2 => n737, A => n278, ZN => n4112);
   U482 : OAI21_X1 port map( B1 => n266, B2 => n738, A => n278, ZN => n4111);
   U483 : OAI21_X1 port map( B1 => n268, B2 => n739, A => n278, ZN => n4110);
   U484 : OAI21_X1 port map( B1 => n266, B2 => n740, A => n278, ZN => n4109);
   U485 : OAI21_X1 port map( B1 => n266, B2 => n741, A => n278, ZN => n4108);
   U486 : OAI21_X1 port map( B1 => n267, B2 => n742, A => n278, ZN => n4107);
   U487 : OAI21_X1 port map( B1 => n267, B2 => n743, A => n278, ZN => n4106);
   U488 : OAI21_X1 port map( B1 => n266, B2 => n744, A => n278, ZN => n4105);
   U489 : OAI21_X1 port map( B1 => n267, B2 => n745, A => n278, ZN => n4104);
   U490 : OAI21_X1 port map( B1 => n267, B2 => n746, A => n278, ZN => n4103);
   U491 : OAI21_X1 port map( B1 => n747, B2 => n748, A => n260, ZN => n715);
   U492 : MUX2_X1 port map( A => n749, B => n281, S => n287, Z => n4102);
   U493 : MUX2_X1 port map( A => n752, B => n288, S => n287, Z => n4101);
   U494 : MUX2_X1 port map( A => n754, B => n291, S => n287, Z => n4100);
   U495 : MUX2_X1 port map( A => n756, B => n294, S => n287, Z => n4099);
   U496 : MUX2_X1 port map( A => n758, B => n297, S => n287, Z => n4098);
   U497 : MUX2_X1 port map( A => n760, B => n300, S => n287, Z => n4097);
   U498 : MUX2_X1 port map( A => n762, B => n303, S => n287, Z => n4096);
   U499 : MUX2_X1 port map( A => n764, B => n306, S => n287, Z => n4095);
   U500 : MUX2_X1 port map( A => n766, B => n309, S => n286, Z => n4094);
   U501 : MUX2_X1 port map( A => n768, B => n312, S => n286, Z => n4093);
   U502 : MUX2_X1 port map( A => n770, B => n315, S => n286, Z => n4092);
   U503 : MUX2_X1 port map( A => n772, B => n318, S => n286, Z => n4091);
   U504 : MUX2_X1 port map( A => n774, B => n321, S => n286, Z => n4090);
   U505 : MUX2_X1 port map( A => n776, B => n324, S => n286, Z => n4089);
   U506 : MUX2_X1 port map( A => n778, B => n327, S => n286, Z => n4088);
   U507 : MUX2_X1 port map( A => n780, B => n330, S => n286, Z => n4087);
   U508 : MUX2_X1 port map( A => n782, B => n333, S => n286, Z => n4086);
   U509 : MUX2_X1 port map( A => n784, B => n336, S => n286, Z => n4085);
   U510 : MUX2_X1 port map( A => n786, B => n339, S => n286, Z => n4084);
   U511 : MUX2_X1 port map( A => n788, B => n342, S => n286, Z => n4083);
   U512 : MUX2_X1 port map( A => n790, B => n345, S => n285, Z => n4082);
   U513 : MUX2_X1 port map( A => n792, B => n348, S => n285, Z => n4081);
   U514 : MUX2_X1 port map( A => n794, B => n351, S => n285, Z => n4080);
   U515 : MUX2_X1 port map( A => n796, B => n354, S => n285, Z => n4079);
   U516 : MUX2_X1 port map( A => n798, B => n357, S => n285, Z => n4078);
   U517 : MUX2_X1 port map( A => n800, B => n360, S => n285, Z => n4077);
   U518 : MUX2_X1 port map( A => n802, B => n363, S => n285, Z => n4076);
   U519 : MUX2_X1 port map( A => n804, B => n366, S => n285, Z => n4075);
   U520 : MUX2_X1 port map( A => n806, B => n369, S => n285, Z => n4074);
   U521 : MUX2_X1 port map( A => n808, B => n372, S => n285, Z => n4073);
   U522 : MUX2_X1 port map( A => n810, B => n375, S => n285, Z => n4072);
   U523 : MUX2_X1 port map( A => n812, B => n378, S => n285, Z => n4071);
   U524 : OAI21_X1 port map( B1 => n814, B2 => n815, A => n261, ZN => n751);
   U525 : MUX2_X1 port map( A => n816, B => n281, S => n384, Z => n4070);
   U526 : MUX2_X1 port map( A => n818, B => n288, S => n384, Z => n4069);
   U527 : MUX2_X1 port map( A => n819, B => n291, S => n384, Z => n4068);
   U528 : MUX2_X1 port map( A => n820, B => n294, S => n384, Z => n4067);
   U529 : MUX2_X1 port map( A => n821, B => n297, S => n384, Z => n4066);
   U530 : MUX2_X1 port map( A => n822, B => n300, S => n384, Z => n4065);
   U531 : MUX2_X1 port map( A => n823, B => n303, S => n384, Z => n4064);
   U532 : MUX2_X1 port map( A => n824, B => n306, S => n384, Z => n4063);
   U533 : MUX2_X1 port map( A => n825, B => n309, S => n383, Z => n4062);
   U534 : MUX2_X1 port map( A => n826, B => n312, S => n383, Z => n4061);
   U535 : MUX2_X1 port map( A => n827, B => n315, S => n383, Z => n4060);
   U536 : MUX2_X1 port map( A => n828, B => n318, S => n383, Z => n4059);
   U537 : MUX2_X1 port map( A => n829, B => n321, S => n383, Z => n4058);
   U538 : MUX2_X1 port map( A => n830, B => n324, S => n383, Z => n4057);
   U539 : MUX2_X1 port map( A => n831, B => n327, S => n383, Z => n4056);
   U540 : MUX2_X1 port map( A => n832, B => n330, S => n383, Z => n4055);
   U541 : MUX2_X1 port map( A => n833, B => n333, S => n383, Z => n4054);
   U542 : MUX2_X1 port map( A => n834, B => n336, S => n383, Z => n4053);
   U543 : MUX2_X1 port map( A => n835, B => n339, S => n383, Z => n4052);
   U544 : MUX2_X1 port map( A => n836, B => n342, S => n383, Z => n4051);
   U545 : MUX2_X1 port map( A => n837, B => n345, S => n382, Z => n4050);
   U546 : MUX2_X1 port map( A => n838, B => n348, S => n382, Z => n4049);
   U547 : MUX2_X1 port map( A => n839, B => n351, S => n382, Z => n4048);
   U548 : MUX2_X1 port map( A => n840, B => n354, S => n382, Z => n4047);
   U549 : MUX2_X1 port map( A => n841, B => n357, S => n382, Z => n4046);
   U550 : MUX2_X1 port map( A => n842, B => n360, S => n382, Z => n4045);
   U551 : MUX2_X1 port map( A => n843, B => n363, S => n382, Z => n4044);
   U552 : MUX2_X1 port map( A => n844, B => n366, S => n382, Z => n4043);
   U553 : MUX2_X1 port map( A => n845, B => n369, S => n382, Z => n4042);
   U554 : MUX2_X1 port map( A => n846, B => n372, S => n382, Z => n4041);
   U555 : MUX2_X1 port map( A => n847, B => n375, S => n382, Z => n4040);
   U556 : MUX2_X1 port map( A => n848, B => n378, S => n382, Z => n4039);
   U557 : OAI21_X1 port map( B1 => n814, B2 => n849, A => n260, ZN => n817);
   U558 : MUX2_X1 port map( A => n5299, B => n281, S => n388, Z => n4038);
   U559 : MUX2_X1 port map( A => n5298, B => n288, S => n388, Z => n4037);
   U560 : MUX2_X1 port map( A => n5297, B => n291, S => n388, Z => n4036);
   U561 : MUX2_X1 port map( A => n5296, B => n294, S => n388, Z => n4035);
   U562 : MUX2_X1 port map( A => n5295, B => n297, S => n388, Z => n4034);
   U563 : MUX2_X1 port map( A => n5294, B => n300, S => n388, Z => n4033);
   U564 : MUX2_X1 port map( A => n5293, B => n303, S => n388, Z => n4032);
   U565 : MUX2_X1 port map( A => n5292, B => n306, S => n388, Z => n4031);
   U566 : MUX2_X1 port map( A => n5291, B => n309, S => n387, Z => n4030);
   U567 : MUX2_X1 port map( A => n5290, B => n312, S => n387, Z => n4029);
   U568 : MUX2_X1 port map( A => n5289, B => n315, S => n387, Z => n4028);
   U569 : MUX2_X1 port map( A => n5288, B => n318, S => n387, Z => n4027);
   U570 : MUX2_X1 port map( A => n5287, B => n321, S => n387, Z => n4026);
   U571 : MUX2_X1 port map( A => n5286, B => n324, S => n387, Z => n4025);
   U572 : MUX2_X1 port map( A => n5285, B => n327, S => n387, Z => n4024);
   U573 : MUX2_X1 port map( A => n5284, B => n330, S => n387, Z => n4023);
   U574 : MUX2_X1 port map( A => n5283, B => n333, S => n387, Z => n4022);
   U575 : MUX2_X1 port map( A => n5282, B => n336, S => n387, Z => n4021);
   U576 : MUX2_X1 port map( A => n5281, B => n339, S => n387, Z => n4020);
   U577 : MUX2_X1 port map( A => n5280, B => n342, S => n387, Z => n4019);
   U578 : MUX2_X1 port map( A => n5279, B => n345, S => n386, Z => n4018);
   U579 : MUX2_X1 port map( A => n5278, B => n348, S => n386, Z => n4017);
   U580 : MUX2_X1 port map( A => n5277, B => n351, S => n386, Z => n4016);
   U581 : MUX2_X1 port map( A => n5276, B => n354, S => n386, Z => n4015);
   U582 : MUX2_X1 port map( A => n5275, B => n357, S => n386, Z => n4014);
   U583 : MUX2_X1 port map( A => n5274, B => n360, S => n386, Z => n4013);
   U584 : MUX2_X1 port map( A => n5273, B => n363, S => n386, Z => n4012);
   U585 : MUX2_X1 port map( A => n5272, B => n366, S => n386, Z => n4011);
   U586 : MUX2_X1 port map( A => n5271, B => n369, S => n386, Z => n4010);
   U587 : MUX2_X1 port map( A => n5270, B => n372, S => n386, Z => n4009);
   U588 : MUX2_X1 port map( A => n5269, B => n375, S => n386, Z => n4008);
   U589 : MUX2_X1 port map( A => n5268, B => n378, S => n386, Z => n4007);
   U590 : OAI21_X1 port map( B1 => n814, B2 => n851, A => n260, ZN => n850);
   U591 : MUX2_X1 port map( A => n5267, B => n281, S => n392, Z => n4006);
   U592 : MUX2_X1 port map( A => n5266, B => n288, S => n392, Z => n4005);
   U593 : MUX2_X1 port map( A => n5265, B => n291, S => n392, Z => n4004);
   U594 : MUX2_X1 port map( A => n5264, B => n294, S => n392, Z => n4003);
   U595 : MUX2_X1 port map( A => n5263, B => n297, S => n392, Z => n4002);
   U596 : MUX2_X1 port map( A => n5262, B => n300, S => n392, Z => n4001);
   U597 : MUX2_X1 port map( A => n5261, B => n303, S => n392, Z => n4000);
   U598 : MUX2_X1 port map( A => n5260, B => n306, S => n392, Z => n3999);
   U599 : MUX2_X1 port map( A => n5259, B => n309, S => n391, Z => n3998);
   U600 : MUX2_X1 port map( A => n5258, B => n312, S => n391, Z => n3997);
   U601 : MUX2_X1 port map( A => n5257, B => n315, S => n391, Z => n3996);
   U602 : MUX2_X1 port map( A => n5256, B => n318, S => n391, Z => n3995);
   U603 : MUX2_X1 port map( A => n5255, B => n321, S => n391, Z => n3994);
   U604 : MUX2_X1 port map( A => n5254, B => n324, S => n391, Z => n3993);
   U605 : MUX2_X1 port map( A => n5253, B => n327, S => n391, Z => n3992);
   U606 : MUX2_X1 port map( A => n5252, B => n330, S => n391, Z => n3991);
   U607 : MUX2_X1 port map( A => n5251, B => n333, S => n391, Z => n3990);
   U608 : MUX2_X1 port map( A => n5250, B => n336, S => n391, Z => n3989);
   U609 : MUX2_X1 port map( A => n5249, B => n339, S => n391, Z => n3988);
   U610 : MUX2_X1 port map( A => n5248, B => n342, S => n391, Z => n3987);
   U611 : MUX2_X1 port map( A => n5247, B => n345, S => n390, Z => n3986);
   U612 : MUX2_X1 port map( A => n5246, B => n348, S => n390, Z => n3985);
   U613 : MUX2_X1 port map( A => n5245, B => n351, S => n390, Z => n3984);
   U614 : MUX2_X1 port map( A => n5244, B => n354, S => n390, Z => n3983);
   U615 : MUX2_X1 port map( A => n5243, B => n357, S => n390, Z => n3982);
   U616 : MUX2_X1 port map( A => n5242, B => n360, S => n390, Z => n3981);
   U617 : MUX2_X1 port map( A => n5241, B => n363, S => n390, Z => n3980);
   U618 : MUX2_X1 port map( A => n5240, B => n366, S => n390, Z => n3979);
   U619 : MUX2_X1 port map( A => n5239, B => n369, S => n390, Z => n3978);
   U620 : MUX2_X1 port map( A => n5238, B => n372, S => n390, Z => n3977);
   U621 : MUX2_X1 port map( A => n5237, B => n375, S => n390, Z => n3976);
   U622 : MUX2_X1 port map( A => n5236, B => n378, S => n390, Z => n3975);
   U623 : OAI21_X1 port map( B1 => n814, B2 => n853, A => n261, ZN => n852);
   U624 : NAND3_X1 port map( A1 => n854, A2 => n855, A3 => n856, ZN => n814);
   U625 : MUX2_X1 port map( A => n857, B => n281, S => n396, Z => n3974);
   U626 : MUX2_X1 port map( A => n859, B => n288, S => n396, Z => n3973);
   U627 : MUX2_X1 port map( A => n860, B => n291, S => n396, Z => n3972);
   U628 : MUX2_X1 port map( A => n861, B => n294, S => n396, Z => n3971);
   U629 : MUX2_X1 port map( A => n862, B => n297, S => n396, Z => n3970);
   U630 : MUX2_X1 port map( A => n863, B => n300, S => n396, Z => n3969);
   U631 : MUX2_X1 port map( A => n864, B => n303, S => n396, Z => n3968);
   U632 : MUX2_X1 port map( A => n865, B => n306, S => n396, Z => n3967);
   U633 : MUX2_X1 port map( A => n866, B => n309, S => n395, Z => n3966);
   U634 : MUX2_X1 port map( A => n867, B => n312, S => n395, Z => n3965);
   U635 : MUX2_X1 port map( A => n868, B => n315, S => n395, Z => n3964);
   U636 : MUX2_X1 port map( A => n869, B => n318, S => n395, Z => n3963);
   U637 : MUX2_X1 port map( A => n870, B => n321, S => n395, Z => n3962);
   U638 : MUX2_X1 port map( A => n871, B => n324, S => n395, Z => n3961);
   U639 : MUX2_X1 port map( A => n872, B => n327, S => n395, Z => n3960);
   U640 : MUX2_X1 port map( A => n873, B => n330, S => n395, Z => n3959);
   U641 : MUX2_X1 port map( A => n874, B => n333, S => n395, Z => n3958);
   U642 : MUX2_X1 port map( A => n875, B => n336, S => n395, Z => n3957);
   U643 : MUX2_X1 port map( A => n876, B => n339, S => n395, Z => n3956);
   U644 : MUX2_X1 port map( A => n877, B => n342, S => n395, Z => n3955);
   U645 : MUX2_X1 port map( A => n878, B => n345, S => n394, Z => n3954);
   U646 : MUX2_X1 port map( A => n879, B => n348, S => n394, Z => n3953);
   U647 : MUX2_X1 port map( A => n880, B => n351, S => n394, Z => n3952);
   U648 : MUX2_X1 port map( A => n881, B => n354, S => n394, Z => n3951);
   U649 : MUX2_X1 port map( A => n882, B => n357, S => n394, Z => n3950);
   U650 : MUX2_X1 port map( A => n883, B => n360, S => n394, Z => n3949);
   U651 : MUX2_X1 port map( A => n884, B => n363, S => n394, Z => n3948);
   U652 : MUX2_X1 port map( A => n885, B => n366, S => n394, Z => n3947);
   U653 : MUX2_X1 port map( A => n886, B => n369, S => n394, Z => n3946);
   U654 : MUX2_X1 port map( A => n887, B => n372, S => n394, Z => n3945);
   U655 : MUX2_X1 port map( A => n888, B => n375, S => n394, Z => n3944);
   U656 : MUX2_X1 port map( A => n889, B => n378, S => n394, Z => n3943);
   U657 : OAI21_X1 port map( B1 => n815, B2 => n890, A => n261, ZN => n858);
   U658 : MUX2_X1 port map( A => n891, B => n281, S => n400, Z => n3942);
   U659 : MUX2_X1 port map( A => n893, B => n288, S => n400, Z => n3941);
   U660 : MUX2_X1 port map( A => n894, B => n291, S => n400, Z => n3940);
   U661 : MUX2_X1 port map( A => n895, B => n294, S => n400, Z => n3939);
   U662 : MUX2_X1 port map( A => n896, B => n297, S => n400, Z => n3938);
   U663 : MUX2_X1 port map( A => n897, B => n300, S => n400, Z => n3937);
   U664 : MUX2_X1 port map( A => n898, B => n303, S => n400, Z => n3936);
   U665 : MUX2_X1 port map( A => n899, B => n306, S => n400, Z => n3935);
   U666 : MUX2_X1 port map( A => n900, B => n309, S => n399, Z => n3934);
   U667 : MUX2_X1 port map( A => n901, B => n312, S => n399, Z => n3933);
   U668 : MUX2_X1 port map( A => n902, B => n315, S => n399, Z => n3932);
   U669 : MUX2_X1 port map( A => n903, B => n318, S => n399, Z => n3931);
   U670 : MUX2_X1 port map( A => n904, B => n321, S => n399, Z => n3930);
   U671 : MUX2_X1 port map( A => n905, B => n324, S => n399, Z => n3929);
   U672 : MUX2_X1 port map( A => n906, B => n327, S => n399, Z => n3928);
   U673 : MUX2_X1 port map( A => n907, B => n330, S => n399, Z => n3927);
   U674 : MUX2_X1 port map( A => n908, B => n333, S => n399, Z => n3926);
   U675 : MUX2_X1 port map( A => n909, B => n336, S => n399, Z => n3925);
   U676 : MUX2_X1 port map( A => n910, B => n339, S => n399, Z => n3924);
   U677 : MUX2_X1 port map( A => n911, B => n342, S => n399, Z => n3923);
   U678 : MUX2_X1 port map( A => n912, B => n345, S => n398, Z => n3922);
   U679 : MUX2_X1 port map( A => n913, B => n348, S => n398, Z => n3921);
   U680 : MUX2_X1 port map( A => n914, B => n351, S => n398, Z => n3920);
   U681 : MUX2_X1 port map( A => n915, B => n354, S => n398, Z => n3919);
   U682 : MUX2_X1 port map( A => n916, B => n357, S => n398, Z => n3918);
   U683 : MUX2_X1 port map( A => n917, B => n360, S => n398, Z => n3917);
   U684 : MUX2_X1 port map( A => n918, B => n363, S => n398, Z => n3916);
   U685 : MUX2_X1 port map( A => n919, B => n366, S => n398, Z => n3915);
   U686 : MUX2_X1 port map( A => n920, B => n369, S => n398, Z => n3914);
   U687 : MUX2_X1 port map( A => n921, B => n372, S => n398, Z => n3913);
   U688 : MUX2_X1 port map( A => n922, B => n375, S => n398, Z => n3912);
   U689 : MUX2_X1 port map( A => n923, B => n378, S => n398, Z => n3911);
   U690 : OAI21_X1 port map( B1 => n849, B2 => n890, A => n261, ZN => n892);
   U691 : MUX2_X1 port map( A => n5171, B => n281, S => n404, Z => n3910);
   U692 : MUX2_X1 port map( A => n5170, B => n288, S => n404, Z => n3909);
   U693 : MUX2_X1 port map( A => n5169, B => n291, S => n404, Z => n3908);
   U694 : MUX2_X1 port map( A => n5168, B => n294, S => n404, Z => n3907);
   U695 : MUX2_X1 port map( A => n5167, B => n297, S => n404, Z => n3906);
   U696 : MUX2_X1 port map( A => n5166, B => n300, S => n404, Z => n3905);
   U697 : MUX2_X1 port map( A => n5165, B => n303, S => n404, Z => n3904);
   U698 : MUX2_X1 port map( A => n5164, B => n306, S => n404, Z => n3903);
   U699 : MUX2_X1 port map( A => n5163, B => n309, S => n403, Z => n3902);
   U700 : MUX2_X1 port map( A => n5162, B => n312, S => n403, Z => n3901);
   U701 : MUX2_X1 port map( A => n5161, B => n315, S => n403, Z => n3900);
   U702 : MUX2_X1 port map( A => n5160, B => n318, S => n403, Z => n3899);
   U703 : MUX2_X1 port map( A => n5159, B => n321, S => n403, Z => n3898);
   U704 : MUX2_X1 port map( A => n5158, B => n324, S => n403, Z => n3897);
   U705 : MUX2_X1 port map( A => n5157, B => n327, S => n403, Z => n3896);
   U706 : MUX2_X1 port map( A => n5156, B => n330, S => n403, Z => n3895);
   U707 : MUX2_X1 port map( A => n5155, B => n333, S => n403, Z => n3894);
   U708 : MUX2_X1 port map( A => n5154, B => n336, S => n403, Z => n3893);
   U709 : MUX2_X1 port map( A => n5153, B => n339, S => n403, Z => n3892);
   U710 : MUX2_X1 port map( A => n5152, B => n342, S => n403, Z => n3891);
   U711 : MUX2_X1 port map( A => n5151, B => n345, S => n402, Z => n3890);
   U712 : MUX2_X1 port map( A => n5150, B => n348, S => n402, Z => n3889);
   U713 : MUX2_X1 port map( A => n5149, B => n351, S => n402, Z => n3888);
   U714 : MUX2_X1 port map( A => n5148, B => n354, S => n402, Z => n3887);
   U715 : MUX2_X1 port map( A => n5147, B => n357, S => n402, Z => n3886);
   U716 : MUX2_X1 port map( A => n5146, B => n360, S => n402, Z => n3885);
   U717 : MUX2_X1 port map( A => n5145, B => n363, S => n402, Z => n3884);
   U718 : MUX2_X1 port map( A => n5144, B => n366, S => n402, Z => n3883);
   U719 : MUX2_X1 port map( A => n5143, B => n369, S => n402, Z => n3882);
   U720 : MUX2_X1 port map( A => n5142, B => n372, S => n402, Z => n3881);
   U721 : MUX2_X1 port map( A => n5141, B => n375, S => n402, Z => n3880);
   U722 : MUX2_X1 port map( A => n5140, B => n378, S => n402, Z => n3879);
   U723 : OAI21_X1 port map( B1 => n851, B2 => n890, A => n261, ZN => n924);
   U724 : MUX2_X1 port map( A => n5139, B => n281, S => n408, Z => n3878);
   U725 : MUX2_X1 port map( A => n5138, B => n288, S => n408, Z => n3877);
   U726 : MUX2_X1 port map( A => n5137, B => n291, S => n408, Z => n3876);
   U727 : MUX2_X1 port map( A => n5136, B => n294, S => n408, Z => n3875);
   U728 : MUX2_X1 port map( A => n5135, B => n297, S => n408, Z => n3874);
   U729 : MUX2_X1 port map( A => n5134, B => n300, S => n408, Z => n3873);
   U730 : MUX2_X1 port map( A => n5133, B => n303, S => n408, Z => n3872);
   U731 : MUX2_X1 port map( A => n5132, B => n306, S => n408, Z => n3871);
   U732 : MUX2_X1 port map( A => n5131, B => n309, S => n407, Z => n3870);
   U733 : MUX2_X1 port map( A => n5130, B => n312, S => n407, Z => n3869);
   U734 : MUX2_X1 port map( A => n5129, B => n315, S => n407, Z => n3868);
   U735 : MUX2_X1 port map( A => n5128, B => n318, S => n407, Z => n3867);
   U736 : MUX2_X1 port map( A => n5127, B => n321, S => n407, Z => n3866);
   U737 : MUX2_X1 port map( A => n5126, B => n324, S => n407, Z => n3865);
   U738 : MUX2_X1 port map( A => n5125, B => n327, S => n407, Z => n3864);
   U739 : MUX2_X1 port map( A => n5124, B => n330, S => n407, Z => n3863);
   U740 : MUX2_X1 port map( A => n5123, B => n333, S => n407, Z => n3862);
   U741 : MUX2_X1 port map( A => n5122, B => n336, S => n407, Z => n3861);
   U742 : MUX2_X1 port map( A => n5121, B => n339, S => n407, Z => n3860);
   U743 : MUX2_X1 port map( A => n5120, B => n342, S => n407, Z => n3859);
   U744 : MUX2_X1 port map( A => n5119, B => n345, S => n406, Z => n3858);
   U745 : MUX2_X1 port map( A => n5118, B => n348, S => n406, Z => n3857);
   U746 : MUX2_X1 port map( A => n5117, B => n351, S => n406, Z => n3856);
   U747 : MUX2_X1 port map( A => n5116, B => n354, S => n406, Z => n3855);
   U748 : MUX2_X1 port map( A => n5115, B => n357, S => n406, Z => n3854);
   U749 : MUX2_X1 port map( A => n5114, B => n360, S => n406, Z => n3853);
   U750 : MUX2_X1 port map( A => n5113, B => n363, S => n406, Z => n3852);
   U751 : MUX2_X1 port map( A => n5112, B => n366, S => n406, Z => n3851);
   U752 : MUX2_X1 port map( A => n5111, B => n369, S => n406, Z => n3850);
   U753 : MUX2_X1 port map( A => n5110, B => n372, S => n406, Z => n3849);
   U754 : MUX2_X1 port map( A => n5109, B => n375, S => n406, Z => n3848);
   U755 : MUX2_X1 port map( A => n5108, B => n378, S => n406, Z => n3847);
   U756 : OAI21_X1 port map( B1 => n853, B2 => n890, A => n260, ZN => n925);
   U757 : NAND3_X1 port map( A1 => n856, A2 => n855, A3 => ADD_WR(2), ZN => 
                           n890);
   U758 : MUX2_X1 port map( A => n926, B => n281, S => n412, Z => n3846);
   U759 : MUX2_X1 port map( A => n928, B => n288, S => n412, Z => n3845);
   U760 : MUX2_X1 port map( A => n929, B => n291, S => n412, Z => n3844);
   U761 : MUX2_X1 port map( A => n930, B => n294, S => n412, Z => n3843);
   U762 : MUX2_X1 port map( A => n931, B => n297, S => n412, Z => n3842);
   U763 : MUX2_X1 port map( A => n932, B => n300, S => n412, Z => n3841);
   U764 : MUX2_X1 port map( A => n933, B => n303, S => n412, Z => n3840);
   U765 : MUX2_X1 port map( A => n934, B => n306, S => n412, Z => n3839);
   U766 : MUX2_X1 port map( A => n935, B => n309, S => n411, Z => n3838);
   U767 : MUX2_X1 port map( A => n936, B => n312, S => n411, Z => n3837);
   U768 : MUX2_X1 port map( A => n937, B => n315, S => n411, Z => n3836);
   U769 : MUX2_X1 port map( A => n938, B => n318, S => n411, Z => n3835);
   U770 : MUX2_X1 port map( A => n939, B => n321, S => n411, Z => n3834);
   U771 : MUX2_X1 port map( A => n940, B => n324, S => n411, Z => n3833);
   U772 : MUX2_X1 port map( A => n941, B => n327, S => n411, Z => n3832);
   U773 : MUX2_X1 port map( A => n942, B => n330, S => n411, Z => n3831);
   U774 : MUX2_X1 port map( A => n943, B => n333, S => n411, Z => n3830);
   U775 : MUX2_X1 port map( A => n944, B => n336, S => n411, Z => n3829);
   U776 : MUX2_X1 port map( A => n945, B => n339, S => n411, Z => n3828);
   U777 : MUX2_X1 port map( A => n946, B => n342, S => n411, Z => n3827);
   U778 : MUX2_X1 port map( A => n947, B => n345, S => n410, Z => n3826);
   U779 : MUX2_X1 port map( A => n948, B => n348, S => n410, Z => n3825);
   U780 : MUX2_X1 port map( A => n949, B => n351, S => n410, Z => n3824);
   U781 : MUX2_X1 port map( A => n950, B => n354, S => n410, Z => n3823);
   U782 : MUX2_X1 port map( A => n951, B => n357, S => n410, Z => n3822);
   U783 : MUX2_X1 port map( A => n952, B => n360, S => n410, Z => n3821);
   U784 : MUX2_X1 port map( A => n953, B => n363, S => n410, Z => n3820);
   U785 : MUX2_X1 port map( A => n954, B => n366, S => n410, Z => n3819);
   U786 : MUX2_X1 port map( A => n955, B => n369, S => n410, Z => n3818);
   U787 : MUX2_X1 port map( A => n956, B => n372, S => n410, Z => n3817);
   U788 : MUX2_X1 port map( A => n957, B => n375, S => n410, Z => n3816);
   U789 : MUX2_X1 port map( A => n958, B => n378, S => n410, Z => n3815);
   U790 : OAI21_X1 port map( B1 => n815, B2 => n959, A => n261, ZN => n927);
   U791 : MUX2_X1 port map( A => n960, B => n281, S => n416, Z => n3814);
   U792 : MUX2_X1 port map( A => n962, B => n288, S => n416, Z => n3813);
   U793 : MUX2_X1 port map( A => n963, B => n291, S => n416, Z => n3812);
   U794 : MUX2_X1 port map( A => n964, B => n294, S => n416, Z => n3811);
   U795 : MUX2_X1 port map( A => n965, B => n297, S => n416, Z => n3810);
   U796 : MUX2_X1 port map( A => n966, B => n300, S => n416, Z => n3809);
   U797 : MUX2_X1 port map( A => n967, B => n303, S => n416, Z => n3808);
   U798 : MUX2_X1 port map( A => n968, B => n306, S => n416, Z => n3807);
   U799 : MUX2_X1 port map( A => n969, B => n309, S => n415, Z => n3806);
   U800 : MUX2_X1 port map( A => n970, B => n312, S => n415, Z => n3805);
   U801 : MUX2_X1 port map( A => n971, B => n315, S => n415, Z => n3804);
   U802 : MUX2_X1 port map( A => n972, B => n318, S => n415, Z => n3803);
   U803 : MUX2_X1 port map( A => n973, B => n321, S => n415, Z => n3802);
   U804 : MUX2_X1 port map( A => n974, B => n324, S => n415, Z => n3801);
   U805 : MUX2_X1 port map( A => n975, B => n327, S => n415, Z => n3800);
   U806 : MUX2_X1 port map( A => n976, B => n330, S => n415, Z => n3799);
   U807 : MUX2_X1 port map( A => n977, B => n333, S => n415, Z => n3798);
   U808 : MUX2_X1 port map( A => n978, B => n336, S => n415, Z => n3797);
   U809 : MUX2_X1 port map( A => n979, B => n339, S => n415, Z => n3796);
   U810 : MUX2_X1 port map( A => n980, B => n342, S => n415, Z => n3795);
   U811 : MUX2_X1 port map( A => n981, B => n345, S => n414, Z => n3794);
   U812 : MUX2_X1 port map( A => n982, B => n348, S => n414, Z => n3793);
   U813 : MUX2_X1 port map( A => n983, B => n351, S => n414, Z => n3792);
   U814 : MUX2_X1 port map( A => n984, B => n354, S => n414, Z => n3791);
   U815 : MUX2_X1 port map( A => n985, B => n357, S => n414, Z => n3790);
   U816 : MUX2_X1 port map( A => n986, B => n360, S => n414, Z => n3789);
   U817 : MUX2_X1 port map( A => n987, B => n363, S => n414, Z => n3788);
   U818 : MUX2_X1 port map( A => n988, B => n366, S => n414, Z => n3787);
   U819 : MUX2_X1 port map( A => n989, B => n369, S => n414, Z => n3786);
   U820 : MUX2_X1 port map( A => n990, B => n372, S => n414, Z => n3785);
   U821 : MUX2_X1 port map( A => n991, B => n375, S => n414, Z => n3784);
   U822 : MUX2_X1 port map( A => n992, B => n378, S => n414, Z => n3783);
   U823 : OAI21_X1 port map( B1 => n849, B2 => n959, A => n261, ZN => n961);
   U824 : MUX2_X1 port map( A => n5043, B => n281, S => n420, Z => n3782);
   U825 : MUX2_X1 port map( A => n5042, B => n288, S => n420, Z => n3781);
   U826 : MUX2_X1 port map( A => n5041, B => n291, S => n420, Z => n3780);
   U827 : MUX2_X1 port map( A => n5040, B => n294, S => n420, Z => n3779);
   U828 : MUX2_X1 port map( A => n5039, B => n297, S => n420, Z => n3778);
   U829 : MUX2_X1 port map( A => n5038, B => n300, S => n420, Z => n3777);
   U830 : MUX2_X1 port map( A => n5037, B => n303, S => n420, Z => n3776);
   U831 : MUX2_X1 port map( A => n5036, B => n306, S => n420, Z => n3775);
   U832 : MUX2_X1 port map( A => n5035, B => n309, S => n419, Z => n3774);
   U833 : MUX2_X1 port map( A => n5034, B => n312, S => n419, Z => n3773);
   U834 : MUX2_X1 port map( A => n5033, B => n315, S => n419, Z => n3772);
   U835 : MUX2_X1 port map( A => n5032, B => n318, S => n419, Z => n3771);
   U836 : MUX2_X1 port map( A => n5031, B => n321, S => n419, Z => n3770);
   U837 : MUX2_X1 port map( A => n5030, B => n324, S => n419, Z => n3769);
   U838 : MUX2_X1 port map( A => n5029, B => n327, S => n419, Z => n3768);
   U839 : MUX2_X1 port map( A => n5028, B => n330, S => n419, Z => n3767);
   U840 : MUX2_X1 port map( A => n5027, B => n333, S => n419, Z => n3766);
   U841 : MUX2_X1 port map( A => n5026, B => n336, S => n419, Z => n3765);
   U842 : MUX2_X1 port map( A => n5025, B => n339, S => n419, Z => n3764);
   U843 : MUX2_X1 port map( A => n5024, B => n342, S => n419, Z => n3763);
   U844 : MUX2_X1 port map( A => n5023, B => n345, S => n418, Z => n3762);
   U845 : MUX2_X1 port map( A => n5022, B => n348, S => n418, Z => n3761);
   U846 : MUX2_X1 port map( A => n5021, B => n351, S => n418, Z => n3760);
   U847 : MUX2_X1 port map( A => n5020, B => n354, S => n418, Z => n3759);
   U848 : MUX2_X1 port map( A => n5019, B => n357, S => n418, Z => n3758);
   U849 : MUX2_X1 port map( A => n5018, B => n360, S => n418, Z => n3757);
   U850 : MUX2_X1 port map( A => n5017, B => n363, S => n418, Z => n3756);
   U851 : MUX2_X1 port map( A => n5016, B => n366, S => n418, Z => n3755);
   U852 : MUX2_X1 port map( A => n5015, B => n369, S => n418, Z => n3754);
   U853 : MUX2_X1 port map( A => n5014, B => n372, S => n418, Z => n3753);
   U854 : MUX2_X1 port map( A => n5013, B => n375, S => n418, Z => n3752);
   U855 : MUX2_X1 port map( A => n5012, B => n378, S => n418, Z => n3751);
   U856 : OAI21_X1 port map( B1 => n851, B2 => n959, A => n260, ZN => n993);
   U857 : MUX2_X1 port map( A => n5011, B => n282, S => n424, Z => n3750);
   U858 : MUX2_X1 port map( A => n5010, B => n289, S => n424, Z => n3749);
   U859 : MUX2_X1 port map( A => n5009, B => n292, S => n424, Z => n3748);
   U860 : MUX2_X1 port map( A => n5008, B => n295, S => n424, Z => n3747);
   U861 : MUX2_X1 port map( A => n5007, B => n298, S => n424, Z => n3746);
   U862 : MUX2_X1 port map( A => n5006, B => n301, S => n424, Z => n3745);
   U863 : MUX2_X1 port map( A => n5005, B => n304, S => n424, Z => n3744);
   U864 : MUX2_X1 port map( A => n5004, B => n307, S => n424, Z => n3743);
   U865 : MUX2_X1 port map( A => n5003, B => n310, S => n423, Z => n3742);
   U866 : MUX2_X1 port map( A => n5002, B => n313, S => n423, Z => n3741);
   U867 : MUX2_X1 port map( A => n5001, B => n316, S => n423, Z => n3740);
   U868 : MUX2_X1 port map( A => n5000, B => n319, S => n423, Z => n3739);
   U869 : MUX2_X1 port map( A => n4999, B => n322, S => n423, Z => n3738);
   U870 : MUX2_X1 port map( A => n4998, B => n325, S => n423, Z => n3737);
   U871 : MUX2_X1 port map( A => n4997, B => n328, S => n423, Z => n3736);
   U872 : MUX2_X1 port map( A => n4996, B => n331, S => n423, Z => n3735);
   U873 : MUX2_X1 port map( A => n4995, B => n334, S => n423, Z => n3734);
   U874 : MUX2_X1 port map( A => n4994, B => n337, S => n423, Z => n3733);
   U875 : MUX2_X1 port map( A => n4993, B => n340, S => n423, Z => n3732);
   U876 : MUX2_X1 port map( A => n4992, B => n343, S => n423, Z => n3731);
   U877 : MUX2_X1 port map( A => n4991, B => n346, S => n422, Z => n3730);
   U878 : MUX2_X1 port map( A => n4990, B => n349, S => n422, Z => n3729);
   U879 : MUX2_X1 port map( A => n4989, B => n352, S => n422, Z => n3728);
   U880 : MUX2_X1 port map( A => n4988, B => n355, S => n422, Z => n3727);
   U881 : MUX2_X1 port map( A => n4987, B => n358, S => n422, Z => n3726);
   U882 : MUX2_X1 port map( A => n4986, B => n361, S => n422, Z => n3725);
   U883 : MUX2_X1 port map( A => n4985, B => n364, S => n422, Z => n3724);
   U884 : MUX2_X1 port map( A => n4984, B => n367, S => n422, Z => n3723);
   U885 : MUX2_X1 port map( A => n4983, B => n370, S => n422, Z => n3722);
   U886 : MUX2_X1 port map( A => n4982, B => n373, S => n422, Z => n3721);
   U887 : MUX2_X1 port map( A => n4981, B => n376, S => n422, Z => n3720);
   U888 : MUX2_X1 port map( A => n4980, B => n379, S => n422, Z => n3719);
   U889 : OAI21_X1 port map( B1 => n853, B2 => n959, A => n261, ZN => n994);
   U890 : NAND3_X1 port map( A1 => n856, A2 => n854, A3 => ADD_WR(3), ZN => 
                           n959);
   U891 : MUX2_X1 port map( A => n995, B => n282, S => n428, Z => n3718);
   U892 : MUX2_X1 port map( A => n997, B => n289, S => n428, Z => n3717);
   U893 : MUX2_X1 port map( A => n998, B => n292, S => n428, Z => n3716);
   U894 : MUX2_X1 port map( A => n999, B => n295, S => n428, Z => n3715);
   U895 : MUX2_X1 port map( A => n1000, B => n298, S => n428, Z => n3714);
   U896 : MUX2_X1 port map( A => n1001, B => n301, S => n428, Z => n3713);
   U897 : MUX2_X1 port map( A => n1002, B => n304, S => n428, Z => n3712);
   U898 : MUX2_X1 port map( A => n1003, B => n307, S => n428, Z => n3711);
   U899 : MUX2_X1 port map( A => n1004, B => n310, S => n427, Z => n3710);
   U900 : MUX2_X1 port map( A => n1005, B => n313, S => n427, Z => n3709);
   U901 : MUX2_X1 port map( A => n1006, B => n316, S => n427, Z => n3708);
   U902 : MUX2_X1 port map( A => n1007, B => n319, S => n427, Z => n3707);
   U903 : MUX2_X1 port map( A => n1008, B => n322, S => n427, Z => n3706);
   U904 : MUX2_X1 port map( A => n1009, B => n325, S => n427, Z => n3705);
   U905 : MUX2_X1 port map( A => n1010, B => n328, S => n427, Z => n3704);
   U906 : MUX2_X1 port map( A => n1011, B => n331, S => n427, Z => n3703);
   U907 : MUX2_X1 port map( A => n1012, B => n334, S => n427, Z => n3702);
   U908 : MUX2_X1 port map( A => n1013, B => n337, S => n427, Z => n3701);
   U909 : MUX2_X1 port map( A => n1014, B => n340, S => n427, Z => n3700);
   U910 : MUX2_X1 port map( A => n1015, B => n343, S => n427, Z => n3699);
   U911 : MUX2_X1 port map( A => n1016, B => n346, S => n426, Z => n3698);
   U912 : MUX2_X1 port map( A => n1017, B => n349, S => n426, Z => n3697);
   U913 : MUX2_X1 port map( A => n1018, B => n352, S => n426, Z => n3696);
   U914 : MUX2_X1 port map( A => n1019, B => n355, S => n426, Z => n3695);
   U915 : MUX2_X1 port map( A => n1020, B => n358, S => n426, Z => n3694);
   U916 : MUX2_X1 port map( A => n1021, B => n361, S => n426, Z => n3693);
   U917 : MUX2_X1 port map( A => n1022, B => n364, S => n426, Z => n3692);
   U918 : MUX2_X1 port map( A => n1023, B => n367, S => n426, Z => n3691);
   U919 : MUX2_X1 port map( A => n1024, B => n370, S => n426, Z => n3690);
   U920 : MUX2_X1 port map( A => n1025, B => n373, S => n426, Z => n3689);
   U921 : MUX2_X1 port map( A => n1026, B => n376, S => n426, Z => n3688);
   U922 : MUX2_X1 port map( A => n1027, B => n379, S => n426, Z => n3687);
   U923 : OAI21_X1 port map( B1 => n815, B2 => n1028, A => n261, ZN => n996);
   U924 : MUX2_X1 port map( A => n1029, B => n282, S => n432, Z => n3686);
   U925 : MUX2_X1 port map( A => n1031, B => n289, S => n432, Z => n3685);
   U926 : MUX2_X1 port map( A => n1032, B => n292, S => n432, Z => n3684);
   U927 : MUX2_X1 port map( A => n1033, B => n295, S => n432, Z => n3683);
   U928 : MUX2_X1 port map( A => n1034, B => n298, S => n432, Z => n3682);
   U929 : MUX2_X1 port map( A => n1035, B => n301, S => n432, Z => n3681);
   U930 : MUX2_X1 port map( A => n1036, B => n304, S => n432, Z => n3680);
   U931 : MUX2_X1 port map( A => n1037, B => n307, S => n432, Z => n3679);
   U932 : MUX2_X1 port map( A => n1038, B => n310, S => n431, Z => n3678);
   U933 : MUX2_X1 port map( A => n1039, B => n313, S => n431, Z => n3677);
   U934 : MUX2_X1 port map( A => n1040, B => n316, S => n431, Z => n3676);
   U935 : MUX2_X1 port map( A => n1041, B => n319, S => n431, Z => n3675);
   U936 : MUX2_X1 port map( A => n1042, B => n322, S => n431, Z => n3674);
   U937 : MUX2_X1 port map( A => n1043, B => n325, S => n431, Z => n3673);
   U938 : MUX2_X1 port map( A => n1044, B => n328, S => n431, Z => n3672);
   U939 : MUX2_X1 port map( A => n1045, B => n331, S => n431, Z => n3671);
   U940 : MUX2_X1 port map( A => n1046, B => n334, S => n431, Z => n3670);
   U941 : MUX2_X1 port map( A => n1047, B => n337, S => n431, Z => n3669);
   U942 : MUX2_X1 port map( A => n1048, B => n340, S => n431, Z => n3668);
   U943 : MUX2_X1 port map( A => n1049, B => n343, S => n431, Z => n3667);
   U944 : MUX2_X1 port map( A => n1050, B => n346, S => n430, Z => n3666);
   U945 : MUX2_X1 port map( A => n1051, B => n349, S => n430, Z => n3665);
   U946 : MUX2_X1 port map( A => n1052, B => n352, S => n430, Z => n3664);
   U947 : MUX2_X1 port map( A => n1053, B => n355, S => n430, Z => n3663);
   U948 : MUX2_X1 port map( A => n1054, B => n358, S => n430, Z => n3662);
   U949 : MUX2_X1 port map( A => n1055, B => n361, S => n430, Z => n3661);
   U950 : MUX2_X1 port map( A => n1056, B => n364, S => n430, Z => n3660);
   U951 : MUX2_X1 port map( A => n1057, B => n367, S => n430, Z => n3659);
   U952 : MUX2_X1 port map( A => n1058, B => n370, S => n430, Z => n3658);
   U953 : MUX2_X1 port map( A => n1059, B => n373, S => n430, Z => n3657);
   U954 : MUX2_X1 port map( A => n1060, B => n376, S => n430, Z => n3656);
   U955 : MUX2_X1 port map( A => n1061, B => n379, S => n430, Z => n3655);
   U956 : OAI21_X1 port map( B1 => n849, B2 => n1028, A => n260, ZN => n1030);
   U957 : MUX2_X1 port map( A => n4915, B => n282, S => n436, Z => n3654);
   U958 : MUX2_X1 port map( A => n4914, B => n289, S => n436, Z => n3653);
   U959 : MUX2_X1 port map( A => n4913, B => n292, S => n436, Z => n3652);
   U960 : MUX2_X1 port map( A => n4912, B => n295, S => n436, Z => n3651);
   U961 : MUX2_X1 port map( A => n4911, B => n298, S => n436, Z => n3650);
   U962 : MUX2_X1 port map( A => n4910, B => n301, S => n436, Z => n3649);
   U963 : MUX2_X1 port map( A => n4909, B => n304, S => n436, Z => n3648);
   U964 : MUX2_X1 port map( A => n4908, B => n307, S => n436, Z => n3647);
   U965 : MUX2_X1 port map( A => n4907, B => n310, S => n435, Z => n3646);
   U966 : MUX2_X1 port map( A => n4906, B => n313, S => n435, Z => n3645);
   U967 : MUX2_X1 port map( A => n4905, B => n316, S => n435, Z => n3644);
   U968 : MUX2_X1 port map( A => n4904, B => n319, S => n435, Z => n3643);
   U969 : MUX2_X1 port map( A => n4903, B => n322, S => n435, Z => n3642);
   U970 : MUX2_X1 port map( A => n4902, B => n325, S => n435, Z => n3641);
   U971 : MUX2_X1 port map( A => n4901, B => n328, S => n435, Z => n3640);
   U972 : MUX2_X1 port map( A => n4900, B => n331, S => n435, Z => n3639);
   U973 : MUX2_X1 port map( A => n4899, B => n334, S => n435, Z => n3638);
   U974 : MUX2_X1 port map( A => n4898, B => n337, S => n435, Z => n3637);
   U975 : MUX2_X1 port map( A => n4897, B => n340, S => n435, Z => n3636);
   U976 : MUX2_X1 port map( A => n4896, B => n343, S => n435, Z => n3635);
   U977 : MUX2_X1 port map( A => n4895, B => n346, S => n434, Z => n3634);
   U978 : MUX2_X1 port map( A => n4894, B => n349, S => n434, Z => n3633);
   U979 : MUX2_X1 port map( A => n4893, B => n352, S => n434, Z => n3632);
   U980 : MUX2_X1 port map( A => n4892, B => n355, S => n434, Z => n3631);
   U981 : MUX2_X1 port map( A => n4891, B => n358, S => n434, Z => n3630);
   U982 : MUX2_X1 port map( A => n4890, B => n361, S => n434, Z => n3629);
   U983 : MUX2_X1 port map( A => n4889, B => n364, S => n434, Z => n3628);
   U984 : MUX2_X1 port map( A => n4888, B => n367, S => n434, Z => n3627);
   U985 : MUX2_X1 port map( A => n4887, B => n370, S => n434, Z => n3626);
   U986 : MUX2_X1 port map( A => n4886, B => n373, S => n434, Z => n3625);
   U987 : MUX2_X1 port map( A => n4885, B => n376, S => n434, Z => n3624);
   U988 : MUX2_X1 port map( A => n4884, B => n379, S => n434, Z => n3623);
   U989 : OAI21_X1 port map( B1 => n851, B2 => n1028, A => n261, ZN => n1062);
   U990 : MUX2_X1 port map( A => n4883, B => n282, S => n440, Z => n3622);
   U991 : MUX2_X1 port map( A => n4882, B => n289, S => n440, Z => n3621);
   U992 : MUX2_X1 port map( A => n4881, B => n292, S => n440, Z => n3620);
   U993 : MUX2_X1 port map( A => n4880, B => n295, S => n440, Z => n3619);
   U994 : MUX2_X1 port map( A => n4879, B => n298, S => n440, Z => n3618);
   U995 : MUX2_X1 port map( A => n4878, B => n301, S => n440, Z => n3617);
   U996 : MUX2_X1 port map( A => n4877, B => n304, S => n440, Z => n3616);
   U997 : MUX2_X1 port map( A => n4876, B => n307, S => n440, Z => n3615);
   U998 : MUX2_X1 port map( A => n4875, B => n310, S => n439, Z => n3614);
   U999 : MUX2_X1 port map( A => n4874, B => n313, S => n439, Z => n3613);
   U1000 : MUX2_X1 port map( A => n4873, B => n316, S => n439, Z => n3612);
   U1001 : MUX2_X1 port map( A => n4872, B => n319, S => n439, Z => n3611);
   U1002 : MUX2_X1 port map( A => n4871, B => n322, S => n439, Z => n3610);
   U1003 : MUX2_X1 port map( A => n4870, B => n325, S => n439, Z => n3609);
   U1004 : MUX2_X1 port map( A => n4869, B => n328, S => n439, Z => n3608);
   U1005 : MUX2_X1 port map( A => n4868, B => n331, S => n439, Z => n3607);
   U1006 : MUX2_X1 port map( A => n4867, B => n334, S => n439, Z => n3606);
   U1007 : MUX2_X1 port map( A => n4866, B => n337, S => n439, Z => n3605);
   U1008 : MUX2_X1 port map( A => n4865, B => n340, S => n439, Z => n3604);
   U1009 : MUX2_X1 port map( A => n4864, B => n343, S => n439, Z => n3603);
   U1010 : MUX2_X1 port map( A => n4863, B => n346, S => n438, Z => n3602);
   U1011 : MUX2_X1 port map( A => n4862, B => n349, S => n438, Z => n3601);
   U1012 : MUX2_X1 port map( A => n4861, B => n352, S => n438, Z => n3600);
   U1013 : MUX2_X1 port map( A => n4860, B => n355, S => n438, Z => n3599);
   U1014 : MUX2_X1 port map( A => n4859, B => n358, S => n438, Z => n3598);
   U1015 : MUX2_X1 port map( A => n4858, B => n361, S => n438, Z => n3597);
   U1016 : MUX2_X1 port map( A => n4857, B => n364, S => n438, Z => n3596);
   U1017 : MUX2_X1 port map( A => n4856, B => n367, S => n438, Z => n3595);
   U1018 : MUX2_X1 port map( A => n4855, B => n370, S => n438, Z => n3594);
   U1019 : MUX2_X1 port map( A => n4854, B => n373, S => n438, Z => n3593);
   U1020 : MUX2_X1 port map( A => n4853, B => n376, S => n438, Z => n3592);
   U1021 : MUX2_X1 port map( A => n4852, B => n379, S => n438, Z => n3591);
   U1022 : OAI21_X1 port map( B1 => n853, B2 => n1028, A => n260, ZN => n1063);
   U1023 : NAND3_X1 port map( A1 => ADD_WR(2), A2 => n856, A3 => ADD_WR(3), ZN 
                           => n1028);
   U1024 : NOR3_X1 port map( A1 => n747, A2 => ADD_WR(4), A3 => n1064, ZN => 
                           n856);
   U1025 : MUX2_X1 port map( A => n1065, B => n282, S => n444, Z => n3590);
   U1026 : MUX2_X1 port map( A => n1067, B => n289, S => n444, Z => n3589);
   U1027 : MUX2_X1 port map( A => n1068, B => n292, S => n444, Z => n3588);
   U1028 : MUX2_X1 port map( A => n1069, B => n295, S => n444, Z => n3587);
   U1029 : MUX2_X1 port map( A => n1070, B => n298, S => n444, Z => n3586);
   U1030 : MUX2_X1 port map( A => n1071, B => n301, S => n444, Z => n3585);
   U1031 : MUX2_X1 port map( A => n1072, B => n304, S => n444, Z => n3584);
   U1032 : MUX2_X1 port map( A => n1073, B => n307, S => n444, Z => n3583);
   U1033 : MUX2_X1 port map( A => n1074, B => n310, S => n443, Z => n3582);
   U1034 : MUX2_X1 port map( A => n1075, B => n313, S => n443, Z => n3581);
   U1035 : MUX2_X1 port map( A => n1076, B => n316, S => n443, Z => n3580);
   U1036 : MUX2_X1 port map( A => n1077, B => n319, S => n443, Z => n3579);
   U1037 : MUX2_X1 port map( A => n1078, B => n322, S => n443, Z => n3578);
   U1038 : MUX2_X1 port map( A => n1079, B => n325, S => n443, Z => n3577);
   U1039 : MUX2_X1 port map( A => n1080, B => n328, S => n443, Z => n3576);
   U1040 : MUX2_X1 port map( A => n1081, B => n331, S => n443, Z => n3575);
   U1041 : MUX2_X1 port map( A => n1082, B => n334, S => n443, Z => n3574);
   U1042 : MUX2_X1 port map( A => n1083, B => n337, S => n443, Z => n3573);
   U1043 : MUX2_X1 port map( A => n1084, B => n340, S => n443, Z => n3572);
   U1044 : MUX2_X1 port map( A => n1085, B => n343, S => n443, Z => n3571);
   U1045 : MUX2_X1 port map( A => n1086, B => n346, S => n442, Z => n3570);
   U1046 : MUX2_X1 port map( A => n1087, B => n349, S => n442, Z => n3569);
   U1047 : MUX2_X1 port map( A => n1088, B => n352, S => n442, Z => n3568);
   U1048 : MUX2_X1 port map( A => n1089, B => n355, S => n442, Z => n3567);
   U1049 : MUX2_X1 port map( A => n1090, B => n358, S => n442, Z => n3566);
   U1050 : MUX2_X1 port map( A => n1091, B => n361, S => n442, Z => n3565);
   U1051 : MUX2_X1 port map( A => n1092, B => n364, S => n442, Z => n3564);
   U1052 : MUX2_X1 port map( A => n1093, B => n367, S => n442, Z => n3563);
   U1053 : MUX2_X1 port map( A => n1094, B => n370, S => n442, Z => n3562);
   U1054 : MUX2_X1 port map( A => n1095, B => n373, S => n442, Z => n3561);
   U1055 : MUX2_X1 port map( A => n1096, B => n376, S => n442, Z => n3560);
   U1056 : MUX2_X1 port map( A => n1097, B => n379, S => n442, Z => n3559);
   U1057 : OAI21_X1 port map( B1 => n815, B2 => n1098, A => n262, ZN => n1066);
   U1058 : MUX2_X1 port map( A => n1099, B => n282, S => n448, Z => n3558);
   U1059 : MUX2_X1 port map( A => n1101, B => n289, S => n448, Z => n3557);
   U1060 : MUX2_X1 port map( A => n1102, B => n292, S => n448, Z => n3556);
   U1061 : MUX2_X1 port map( A => n1103, B => n295, S => n448, Z => n3555);
   U1062 : MUX2_X1 port map( A => n1104, B => n298, S => n448, Z => n3554);
   U1063 : MUX2_X1 port map( A => n1105, B => n301, S => n448, Z => n3553);
   U1064 : MUX2_X1 port map( A => n1106, B => n304, S => n448, Z => n3552);
   U1065 : MUX2_X1 port map( A => n1107, B => n307, S => n448, Z => n3551);
   U1066 : MUX2_X1 port map( A => n1108, B => n310, S => n447, Z => n3550);
   U1067 : MUX2_X1 port map( A => n1109, B => n313, S => n447, Z => n3549);
   U1068 : MUX2_X1 port map( A => n1110, B => n316, S => n447, Z => n3548);
   U1069 : MUX2_X1 port map( A => n1111, B => n319, S => n447, Z => n3547);
   U1070 : MUX2_X1 port map( A => n1112, B => n322, S => n447, Z => n3546);
   U1071 : MUX2_X1 port map( A => n1113, B => n325, S => n447, Z => n3545);
   U1072 : MUX2_X1 port map( A => n1114, B => n328, S => n447, Z => n3544);
   U1073 : MUX2_X1 port map( A => n1115, B => n331, S => n447, Z => n3543);
   U1074 : MUX2_X1 port map( A => n1116, B => n334, S => n447, Z => n3542);
   U1075 : MUX2_X1 port map( A => n1117, B => n337, S => n447, Z => n3541);
   U1076 : MUX2_X1 port map( A => n1118, B => n340, S => n447, Z => n3540);
   U1077 : MUX2_X1 port map( A => n1119, B => n343, S => n447, Z => n3539);
   U1078 : MUX2_X1 port map( A => n1120, B => n346, S => n446, Z => n3538);
   U1079 : MUX2_X1 port map( A => n1121, B => n349, S => n446, Z => n3537);
   U1080 : MUX2_X1 port map( A => n1122, B => n352, S => n446, Z => n3536);
   U1081 : MUX2_X1 port map( A => n1123, B => n355, S => n446, Z => n3535);
   U1082 : MUX2_X1 port map( A => n1124, B => n358, S => n446, Z => n3534);
   U1083 : MUX2_X1 port map( A => n1125, B => n361, S => n446, Z => n3533);
   U1084 : MUX2_X1 port map( A => n1126, B => n364, S => n446, Z => n3532);
   U1085 : MUX2_X1 port map( A => n1127, B => n367, S => n446, Z => n3531);
   U1086 : MUX2_X1 port map( A => n1128, B => n370, S => n446, Z => n3530);
   U1087 : MUX2_X1 port map( A => n1129, B => n373, S => n446, Z => n3529);
   U1088 : MUX2_X1 port map( A => n1130, B => n376, S => n446, Z => n3528);
   U1089 : MUX2_X1 port map( A => n1131, B => n379, S => n446, Z => n3527);
   U1090 : OAI21_X1 port map( B1 => n849, B2 => n1098, A => n262, ZN => n1100);
   U1091 : MUX2_X1 port map( A => n4787, B => n282, S => n452, Z => n3526);
   U1092 : MUX2_X1 port map( A => n4786, B => n289, S => n452, Z => n3525);
   U1093 : MUX2_X1 port map( A => n4785, B => n292, S => n452, Z => n3524);
   U1094 : MUX2_X1 port map( A => n4784, B => n295, S => n452, Z => n3523);
   U1095 : MUX2_X1 port map( A => n4783, B => n298, S => n452, Z => n3522);
   U1096 : MUX2_X1 port map( A => n4782, B => n301, S => n452, Z => n3521);
   U1097 : MUX2_X1 port map( A => n4781, B => n304, S => n452, Z => n3520);
   U1098 : MUX2_X1 port map( A => n4780, B => n307, S => n452, Z => n3519);
   U1099 : MUX2_X1 port map( A => n4779, B => n310, S => n451, Z => n3518);
   U1100 : MUX2_X1 port map( A => n4778, B => n313, S => n451, Z => n3517);
   U1101 : MUX2_X1 port map( A => n4777, B => n316, S => n451, Z => n3516);
   U1102 : MUX2_X1 port map( A => n4776, B => n319, S => n451, Z => n3515);
   U1103 : MUX2_X1 port map( A => n4775, B => n322, S => n451, Z => n3514);
   U1104 : MUX2_X1 port map( A => n4774, B => n325, S => n451, Z => n3513);
   U1105 : MUX2_X1 port map( A => n4773, B => n328, S => n451, Z => n3512);
   U1106 : MUX2_X1 port map( A => n4772, B => n331, S => n451, Z => n3511);
   U1107 : MUX2_X1 port map( A => n4771, B => n334, S => n451, Z => n3510);
   U1108 : MUX2_X1 port map( A => n4770, B => n337, S => n451, Z => n3509);
   U1109 : MUX2_X1 port map( A => n4769, B => n340, S => n451, Z => n3508);
   U1110 : MUX2_X1 port map( A => n4768, B => n343, S => n451, Z => n3507);
   U1111 : MUX2_X1 port map( A => n4767, B => n346, S => n450, Z => n3506);
   U1112 : MUX2_X1 port map( A => n4766, B => n349, S => n450, Z => n3505);
   U1113 : MUX2_X1 port map( A => n4765, B => n352, S => n450, Z => n3504);
   U1114 : MUX2_X1 port map( A => n4764, B => n355, S => n450, Z => n3503);
   U1115 : MUX2_X1 port map( A => n4763, B => n358, S => n450, Z => n3502);
   U1116 : MUX2_X1 port map( A => n4762, B => n361, S => n450, Z => n3501);
   U1117 : MUX2_X1 port map( A => n4761, B => n364, S => n450, Z => n3500);
   U1118 : MUX2_X1 port map( A => n4760, B => n367, S => n450, Z => n3499);
   U1119 : MUX2_X1 port map( A => n4759, B => n370, S => n450, Z => n3498);
   U1120 : MUX2_X1 port map( A => n4758, B => n373, S => n450, Z => n3497);
   U1121 : MUX2_X1 port map( A => n4757, B => n376, S => n450, Z => n3496);
   U1122 : MUX2_X1 port map( A => n4756, B => n379, S => n450, Z => n3495);
   U1123 : OAI21_X1 port map( B1 => n851, B2 => n1098, A => n260, ZN => n1132);
   U1124 : MUX2_X1 port map( A => n4755, B => n282, S => n456, Z => n3494);
   U1125 : MUX2_X1 port map( A => n4754, B => n289, S => n456, Z => n3493);
   U1126 : MUX2_X1 port map( A => n4753, B => n292, S => n456, Z => n3492);
   U1127 : MUX2_X1 port map( A => n4752, B => n295, S => n456, Z => n3491);
   U1128 : MUX2_X1 port map( A => n4751, B => n298, S => n456, Z => n3490);
   U1129 : MUX2_X1 port map( A => n4750, B => n301, S => n456, Z => n3489);
   U1130 : MUX2_X1 port map( A => n4749, B => n304, S => n456, Z => n3488);
   U1131 : MUX2_X1 port map( A => n4748, B => n307, S => n456, Z => n3487);
   U1132 : MUX2_X1 port map( A => n4747, B => n310, S => n455, Z => n3486);
   U1133 : MUX2_X1 port map( A => n4746, B => n313, S => n455, Z => n3485);
   U1134 : MUX2_X1 port map( A => n4745, B => n316, S => n455, Z => n3484);
   U1135 : MUX2_X1 port map( A => n4744, B => n319, S => n455, Z => n3483);
   U1136 : MUX2_X1 port map( A => n4743, B => n322, S => n455, Z => n3482);
   U1137 : MUX2_X1 port map( A => n4742, B => n325, S => n455, Z => n3481);
   U1138 : MUX2_X1 port map( A => n4741, B => n328, S => n455, Z => n3480);
   U1139 : MUX2_X1 port map( A => n4740, B => n331, S => n455, Z => n3479);
   U1140 : MUX2_X1 port map( A => n4739, B => n334, S => n455, Z => n3478);
   U1141 : MUX2_X1 port map( A => n4738, B => n337, S => n455, Z => n3477);
   U1142 : MUX2_X1 port map( A => n4737, B => n340, S => n455, Z => n3476);
   U1143 : MUX2_X1 port map( A => n4736, B => n343, S => n455, Z => n3475);
   U1144 : MUX2_X1 port map( A => n4735, B => n346, S => n454, Z => n3474);
   U1145 : MUX2_X1 port map( A => n4734, B => n349, S => n454, Z => n3473);
   U1146 : MUX2_X1 port map( A => n4733, B => n352, S => n454, Z => n3472);
   U1147 : MUX2_X1 port map( A => n4732, B => n355, S => n454, Z => n3471);
   U1148 : MUX2_X1 port map( A => n4731, B => n358, S => n454, Z => n3470);
   U1149 : MUX2_X1 port map( A => n4730, B => n361, S => n454, Z => n3469);
   U1150 : MUX2_X1 port map( A => n4729, B => n364, S => n454, Z => n3468);
   U1151 : MUX2_X1 port map( A => n4728, B => n367, S => n454, Z => n3467);
   U1152 : MUX2_X1 port map( A => n4727, B => n370, S => n454, Z => n3466);
   U1153 : MUX2_X1 port map( A => n4726, B => n373, S => n454, Z => n3465);
   U1154 : MUX2_X1 port map( A => n4725, B => n376, S => n454, Z => n3464);
   U1155 : MUX2_X1 port map( A => n4724, B => n379, S => n454, Z => n3463);
   U1156 : OAI21_X1 port map( B1 => n853, B2 => n1098, A => n261, ZN => n1133);
   U1157 : NAND3_X1 port map( A1 => n854, A2 => n855, A3 => n1134, ZN => n1098)
                           ;
   U1158 : MUX2_X1 port map( A => n1135, B => n282, S => n460, Z => n3462);
   U1159 : MUX2_X1 port map( A => n1137, B => n289, S => n460, Z => n3461);
   U1160 : MUX2_X1 port map( A => n1138, B => n292, S => n460, Z => n3460);
   U1161 : MUX2_X1 port map( A => n1139, B => n295, S => n460, Z => n3459);
   U1162 : MUX2_X1 port map( A => n1140, B => n298, S => n460, Z => n3458);
   U1163 : MUX2_X1 port map( A => n1141, B => n301, S => n460, Z => n3457);
   U1164 : MUX2_X1 port map( A => n1142, B => n304, S => n460, Z => n3456);
   U1165 : MUX2_X1 port map( A => n1143, B => n307, S => n460, Z => n3455);
   U1166 : MUX2_X1 port map( A => n1144, B => n310, S => n459, Z => n3454);
   U1167 : MUX2_X1 port map( A => n1145, B => n313, S => n459, Z => n3453);
   U1168 : MUX2_X1 port map( A => n1146, B => n316, S => n459, Z => n3452);
   U1169 : MUX2_X1 port map( A => n1147, B => n319, S => n459, Z => n3451);
   U1170 : MUX2_X1 port map( A => n1148, B => n322, S => n459, Z => n3450);
   U1171 : MUX2_X1 port map( A => n1149, B => n325, S => n459, Z => n3449);
   U1172 : MUX2_X1 port map( A => n1150, B => n328, S => n459, Z => n3448);
   U1173 : MUX2_X1 port map( A => n1151, B => n331, S => n459, Z => n3447);
   U1174 : MUX2_X1 port map( A => n1152, B => n334, S => n459, Z => n3446);
   U1175 : MUX2_X1 port map( A => n1153, B => n337, S => n459, Z => n3445);
   U1176 : MUX2_X1 port map( A => n1154, B => n340, S => n459, Z => n3444);
   U1177 : MUX2_X1 port map( A => n1155, B => n343, S => n459, Z => n3443);
   U1178 : MUX2_X1 port map( A => n1156, B => n346, S => n458, Z => n3442);
   U1179 : MUX2_X1 port map( A => n1157, B => n349, S => n458, Z => n3441);
   U1180 : MUX2_X1 port map( A => n1158, B => n352, S => n458, Z => n3440);
   U1181 : MUX2_X1 port map( A => n1159, B => n355, S => n458, Z => n3439);
   U1182 : MUX2_X1 port map( A => n1160, B => n358, S => n458, Z => n3438);
   U1183 : MUX2_X1 port map( A => n1161, B => n361, S => n458, Z => n3437);
   U1184 : MUX2_X1 port map( A => n1162, B => n364, S => n458, Z => n3436);
   U1185 : MUX2_X1 port map( A => n1163, B => n367, S => n458, Z => n3435);
   U1186 : MUX2_X1 port map( A => n1164, B => n370, S => n458, Z => n3434);
   U1187 : MUX2_X1 port map( A => n1165, B => n373, S => n458, Z => n3433);
   U1188 : MUX2_X1 port map( A => n1166, B => n376, S => n458, Z => n3432);
   U1189 : MUX2_X1 port map( A => n1167, B => n379, S => n458, Z => n3431);
   U1190 : OAI21_X1 port map( B1 => n815, B2 => n1168, A => n262, ZN => n1136);
   U1191 : MUX2_X1 port map( A => n1169, B => n282, S => n464, Z => n3430);
   U1192 : MUX2_X1 port map( A => n1171, B => n289, S => n464, Z => n3429);
   U1193 : MUX2_X1 port map( A => n1172, B => n292, S => n464, Z => n3428);
   U1194 : MUX2_X1 port map( A => n1173, B => n295, S => n464, Z => n3427);
   U1195 : MUX2_X1 port map( A => n1174, B => n298, S => n464, Z => n3426);
   U1196 : MUX2_X1 port map( A => n1175, B => n301, S => n464, Z => n3425);
   U1197 : MUX2_X1 port map( A => n1176, B => n304, S => n464, Z => n3424);
   U1198 : MUX2_X1 port map( A => n1177, B => n307, S => n464, Z => n3423);
   U1199 : MUX2_X1 port map( A => n1178, B => n310, S => n463, Z => n3422);
   U1200 : MUX2_X1 port map( A => n1179, B => n313, S => n463, Z => n3421);
   U1201 : MUX2_X1 port map( A => n1180, B => n316, S => n463, Z => n3420);
   U1202 : MUX2_X1 port map( A => n1181, B => n319, S => n463, Z => n3419);
   U1203 : MUX2_X1 port map( A => n1182, B => n322, S => n463, Z => n3418);
   U1204 : MUX2_X1 port map( A => n1183, B => n325, S => n463, Z => n3417);
   U1205 : MUX2_X1 port map( A => n1184, B => n328, S => n463, Z => n3416);
   U1206 : MUX2_X1 port map( A => n1185, B => n331, S => n463, Z => n3415);
   U1207 : MUX2_X1 port map( A => n1186, B => n334, S => n463, Z => n3414);
   U1208 : MUX2_X1 port map( A => n1187, B => n337, S => n463, Z => n3413);
   U1209 : MUX2_X1 port map( A => n1188, B => n340, S => n463, Z => n3412);
   U1210 : MUX2_X1 port map( A => n1189, B => n343, S => n463, Z => n3411);
   U1211 : MUX2_X1 port map( A => n1190, B => n346, S => n462, Z => n3410);
   U1212 : MUX2_X1 port map( A => n1191, B => n349, S => n462, Z => n3409);
   U1213 : MUX2_X1 port map( A => n1192, B => n352, S => n462, Z => n3408);
   U1214 : MUX2_X1 port map( A => n1193, B => n355, S => n462, Z => n3407);
   U1215 : MUX2_X1 port map( A => n1194, B => n358, S => n462, Z => n3406);
   U1216 : MUX2_X1 port map( A => n1195, B => n361, S => n462, Z => n3405);
   U1217 : MUX2_X1 port map( A => n1196, B => n364, S => n462, Z => n3404);
   U1218 : MUX2_X1 port map( A => n1197, B => n367, S => n462, Z => n3403);
   U1219 : MUX2_X1 port map( A => n1198, B => n370, S => n462, Z => n3402);
   U1220 : MUX2_X1 port map( A => n1199, B => n373, S => n462, Z => n3401);
   U1221 : MUX2_X1 port map( A => n1200, B => n376, S => n462, Z => n3400);
   U1222 : MUX2_X1 port map( A => n1201, B => n379, S => n462, Z => n3399);
   U1223 : OAI21_X1 port map( B1 => n849, B2 => n1168, A => n262, ZN => n1170);
   U1224 : MUX2_X1 port map( A => n4659, B => n283, S => n468, Z => n3398);
   U1225 : MUX2_X1 port map( A => n4658, B => n290, S => n468, Z => n3397);
   U1226 : MUX2_X1 port map( A => n4657, B => n293, S => n468, Z => n3396);
   U1227 : MUX2_X1 port map( A => n4656, B => n296, S => n468, Z => n3395);
   U1228 : MUX2_X1 port map( A => n4655, B => n299, S => n468, Z => n3394);
   U1229 : MUX2_X1 port map( A => n4654, B => n302, S => n468, Z => n3393);
   U1230 : MUX2_X1 port map( A => n4653, B => n305, S => n468, Z => n3392);
   U1231 : MUX2_X1 port map( A => n4652, B => n308, S => n468, Z => n3391);
   U1232 : MUX2_X1 port map( A => n4651, B => n311, S => n467, Z => n3390);
   U1233 : MUX2_X1 port map( A => n4650, B => n314, S => n467, Z => n3389);
   U1234 : MUX2_X1 port map( A => n4649, B => n317, S => n467, Z => n3388);
   U1235 : MUX2_X1 port map( A => n4648, B => n320, S => n467, Z => n3387);
   U1236 : MUX2_X1 port map( A => n4647, B => n323, S => n467, Z => n3386);
   U1237 : MUX2_X1 port map( A => n4646, B => n326, S => n467, Z => n3385);
   U1238 : MUX2_X1 port map( A => n4645, B => n329, S => n467, Z => n3384);
   U1239 : MUX2_X1 port map( A => n4644, B => n332, S => n467, Z => n3383);
   U1240 : MUX2_X1 port map( A => n4643, B => n335, S => n467, Z => n3382);
   U1241 : MUX2_X1 port map( A => n4642, B => n338, S => n467, Z => n3381);
   U1242 : MUX2_X1 port map( A => n4641, B => n341, S => n467, Z => n3380);
   U1243 : MUX2_X1 port map( A => n4640, B => n344, S => n467, Z => n3379);
   U1244 : MUX2_X1 port map( A => n4639, B => n347, S => n466, Z => n3378);
   U1245 : MUX2_X1 port map( A => n4638, B => n350, S => n466, Z => n3377);
   U1246 : MUX2_X1 port map( A => n4637, B => n353, S => n466, Z => n3376);
   U1247 : MUX2_X1 port map( A => n4636, B => n356, S => n466, Z => n3375);
   U1248 : MUX2_X1 port map( A => n4635, B => n359, S => n466, Z => n3374);
   U1249 : MUX2_X1 port map( A => n4634, B => n362, S => n466, Z => n3373);
   U1250 : MUX2_X1 port map( A => n4633, B => n365, S => n466, Z => n3372);
   U1251 : MUX2_X1 port map( A => n4632, B => n368, S => n466, Z => n3371);
   U1252 : MUX2_X1 port map( A => n4631, B => n371, S => n466, Z => n3370);
   U1253 : MUX2_X1 port map( A => n4630, B => n374, S => n466, Z => n3369);
   U1254 : MUX2_X1 port map( A => n4629, B => n377, S => n466, Z => n3368);
   U1255 : MUX2_X1 port map( A => n4628, B => n380, S => n466, Z => n3367);
   U1256 : OAI21_X1 port map( B1 => n851, B2 => n1168, A => n262, ZN => n1202);
   U1257 : MUX2_X1 port map( A => n4627, B => n283, S => n472, Z => n3366);
   U1258 : MUX2_X1 port map( A => n4626, B => n290, S => n472, Z => n3365);
   U1259 : MUX2_X1 port map( A => n4625, B => n293, S => n472, Z => n3364);
   U1260 : MUX2_X1 port map( A => n4624, B => n296, S => n472, Z => n3363);
   U1261 : MUX2_X1 port map( A => n4623, B => n299, S => n472, Z => n3362);
   U1262 : MUX2_X1 port map( A => n4622, B => n302, S => n472, Z => n3361);
   U1263 : MUX2_X1 port map( A => n4621, B => n305, S => n472, Z => n3360);
   U1264 : MUX2_X1 port map( A => n4620, B => n308, S => n472, Z => n3359);
   U1265 : MUX2_X1 port map( A => n4619, B => n311, S => n471, Z => n3358);
   U1266 : MUX2_X1 port map( A => n4618, B => n314, S => n471, Z => n3357);
   U1267 : MUX2_X1 port map( A => n4617, B => n317, S => n471, Z => n3356);
   U1268 : MUX2_X1 port map( A => n4616, B => n320, S => n471, Z => n3355);
   U1269 : MUX2_X1 port map( A => n4615, B => n323, S => n471, Z => n3354);
   U1270 : MUX2_X1 port map( A => n4614, B => n326, S => n471, Z => n3353);
   U1271 : MUX2_X1 port map( A => n4613, B => n329, S => n471, Z => n3352);
   U1272 : MUX2_X1 port map( A => n4612, B => n332, S => n471, Z => n3351);
   U1273 : MUX2_X1 port map( A => n4611, B => n335, S => n471, Z => n3350);
   U1274 : MUX2_X1 port map( A => n4610, B => n338, S => n471, Z => n3349);
   U1275 : MUX2_X1 port map( A => n4609, B => n341, S => n471, Z => n3348);
   U1276 : MUX2_X1 port map( A => n4608, B => n344, S => n471, Z => n3347);
   U1277 : MUX2_X1 port map( A => n4607, B => n347, S => n470, Z => n3346);
   U1278 : MUX2_X1 port map( A => n4606, B => n350, S => n470, Z => n3345);
   U1279 : MUX2_X1 port map( A => n4605, B => n353, S => n470, Z => n3344);
   U1280 : MUX2_X1 port map( A => n4604, B => n356, S => n470, Z => n3343);
   U1281 : MUX2_X1 port map( A => n4603, B => n359, S => n470, Z => n3342);
   U1282 : MUX2_X1 port map( A => n4602, B => n362, S => n470, Z => n3341);
   U1283 : MUX2_X1 port map( A => n4601, B => n365, S => n470, Z => n3340);
   U1284 : MUX2_X1 port map( A => n4600, B => n368, S => n470, Z => n3339);
   U1285 : MUX2_X1 port map( A => n4599, B => n371, S => n470, Z => n3338);
   U1286 : MUX2_X1 port map( A => n4598, B => n374, S => n470, Z => n3337);
   U1287 : MUX2_X1 port map( A => n4597, B => n377, S => n470, Z => n3336);
   U1288 : MUX2_X1 port map( A => n4596, B => n380, S => n470, Z => n3335);
   U1289 : OAI21_X1 port map( B1 => n853, B2 => n1168, A => n260, ZN => n1203);
   U1290 : NAND3_X1 port map( A1 => ADD_WR(2), A2 => n855, A3 => n1134, ZN => 
                           n1168);
   U1291 : INV_X1 port map( A => ADD_WR(3), ZN => n855);
   U1292 : MUX2_X1 port map( A => n4595, B => n283, S => n476, Z => n3334);
   U1293 : MUX2_X1 port map( A => n4594, B => n290, S => n476, Z => n3333);
   U1294 : MUX2_X1 port map( A => n4593, B => n293, S => n476, Z => n3332);
   U1295 : MUX2_X1 port map( A => n4592, B => n296, S => n476, Z => n3331);
   U1296 : MUX2_X1 port map( A => n4591, B => n299, S => n476, Z => n3330);
   U1297 : MUX2_X1 port map( A => n4590, B => n302, S => n476, Z => n3329);
   U1298 : MUX2_X1 port map( A => n4589, B => n305, S => n476, Z => n3328);
   U1299 : MUX2_X1 port map( A => n4588, B => n308, S => n476, Z => n3327);
   U1300 : MUX2_X1 port map( A => n4587, B => n311, S => n475, Z => n3326);
   U1301 : MUX2_X1 port map( A => n4586, B => n314, S => n475, Z => n3325);
   U1302 : MUX2_X1 port map( A => n4585, B => n317, S => n475, Z => n3324);
   U1303 : MUX2_X1 port map( A => n4584, B => n320, S => n475, Z => n3323);
   U1304 : MUX2_X1 port map( A => n4583, B => n323, S => n475, Z => n3322);
   U1305 : MUX2_X1 port map( A => n4582, B => n326, S => n475, Z => n3321);
   U1306 : MUX2_X1 port map( A => n4581, B => n329, S => n475, Z => n3320);
   U1307 : MUX2_X1 port map( A => n4580, B => n332, S => n475, Z => n3319);
   U1308 : MUX2_X1 port map( A => n4579, B => n335, S => n475, Z => n3318);
   U1309 : MUX2_X1 port map( A => n4578, B => n338, S => n475, Z => n3317);
   U1310 : MUX2_X1 port map( A => n4577, B => n341, S => n475, Z => n3316);
   U1311 : MUX2_X1 port map( A => n4576, B => n344, S => n475, Z => n3315);
   U1312 : MUX2_X1 port map( A => n4575, B => n347, S => n474, Z => n3314);
   U1313 : MUX2_X1 port map( A => n4574, B => n350, S => n474, Z => n3313);
   U1314 : MUX2_X1 port map( A => n4573, B => n353, S => n474, Z => n3312);
   U1315 : MUX2_X1 port map( A => n4572, B => n356, S => n474, Z => n3311);
   U1316 : MUX2_X1 port map( A => n4571, B => n359, S => n474, Z => n3310);
   U1317 : MUX2_X1 port map( A => n4570, B => n362, S => n474, Z => n3309);
   U1318 : MUX2_X1 port map( A => n4569, B => n365, S => n474, Z => n3308);
   U1319 : MUX2_X1 port map( A => n4568, B => n368, S => n474, Z => n3307);
   U1320 : MUX2_X1 port map( A => n4567, B => n371, S => n474, Z => n3306);
   U1321 : MUX2_X1 port map( A => n4566, B => n374, S => n474, Z => n3305);
   U1322 : MUX2_X1 port map( A => n4565, B => n377, S => n474, Z => n3304);
   U1323 : MUX2_X1 port map( A => n4564, B => n380, S => n474, Z => n3303);
   U1324 : OAI21_X1 port map( B1 => n815, B2 => n1205, A => n262, ZN => n1204);
   U1325 : MUX2_X1 port map( A => n4563, B => n283, S => n480, Z => n3302);
   U1326 : MUX2_X1 port map( A => n4562, B => n290, S => n480, Z => n3301);
   U1327 : MUX2_X1 port map( A => n4561, B => n293, S => n480, Z => n3300);
   U1328 : MUX2_X1 port map( A => n4560, B => n296, S => n480, Z => n3299);
   U1329 : MUX2_X1 port map( A => n4559, B => n299, S => n480, Z => n3298);
   U1330 : MUX2_X1 port map( A => n4558, B => n302, S => n480, Z => n3297);
   U1331 : MUX2_X1 port map( A => n4557, B => n305, S => n480, Z => n3296);
   U1332 : MUX2_X1 port map( A => n4556, B => n308, S => n480, Z => n3295);
   U1333 : MUX2_X1 port map( A => n4555, B => n311, S => n479, Z => n3294);
   U1334 : MUX2_X1 port map( A => n4554, B => n314, S => n479, Z => n3293);
   U1335 : MUX2_X1 port map( A => n4553, B => n317, S => n479, Z => n3292);
   U1336 : MUX2_X1 port map( A => n4552, B => n320, S => n479, Z => n3291);
   U1337 : MUX2_X1 port map( A => n4551, B => n323, S => n479, Z => n3290);
   U1338 : MUX2_X1 port map( A => n4550, B => n326, S => n479, Z => n3289);
   U1339 : MUX2_X1 port map( A => n4549, B => n329, S => n479, Z => n3288);
   U1340 : MUX2_X1 port map( A => n4548, B => n332, S => n479, Z => n3287);
   U1341 : MUX2_X1 port map( A => n4547, B => n335, S => n479, Z => n3286);
   U1342 : MUX2_X1 port map( A => n4546, B => n338, S => n479, Z => n3285);
   U1343 : MUX2_X1 port map( A => n4545, B => n341, S => n479, Z => n3284);
   U1344 : MUX2_X1 port map( A => n4544, B => n344, S => n479, Z => n3283);
   U1345 : MUX2_X1 port map( A => n4543, B => n347, S => n478, Z => n3282);
   U1346 : MUX2_X1 port map( A => n4542, B => n350, S => n478, Z => n3281);
   U1347 : MUX2_X1 port map( A => n4541, B => n353, S => n478, Z => n3280);
   U1348 : MUX2_X1 port map( A => n4540, B => n356, S => n478, Z => n3279);
   U1349 : MUX2_X1 port map( A => n4539, B => n359, S => n478, Z => n3278);
   U1350 : MUX2_X1 port map( A => n4538, B => n362, S => n478, Z => n3277);
   U1351 : MUX2_X1 port map( A => n4537, B => n365, S => n478, Z => n3276);
   U1352 : MUX2_X1 port map( A => n4536, B => n368, S => n478, Z => n3275);
   U1353 : MUX2_X1 port map( A => n4535, B => n371, S => n478, Z => n3274);
   U1354 : MUX2_X1 port map( A => n4534, B => n374, S => n478, Z => n3273);
   U1355 : MUX2_X1 port map( A => n4533, B => n377, S => n478, Z => n3272);
   U1356 : MUX2_X1 port map( A => n4532, B => n380, S => n478, Z => n3271);
   U1357 : OAI21_X1 port map( B1 => n849, B2 => n1205, A => n261, ZN => n1206);
   U1358 : MUX2_X1 port map( A => n1207, B => n283, S => n484, Z => n3270);
   U1359 : MUX2_X1 port map( A => n1209, B => n290, S => n484, Z => n3269);
   U1360 : MUX2_X1 port map( A => n1210, B => n293, S => n484, Z => n3268);
   U1361 : MUX2_X1 port map( A => n1211, B => n296, S => n484, Z => n3267);
   U1362 : MUX2_X1 port map( A => n1212, B => n299, S => n484, Z => n3266);
   U1363 : MUX2_X1 port map( A => n1213, B => n302, S => n484, Z => n3265);
   U1364 : MUX2_X1 port map( A => n1214, B => n305, S => n484, Z => n3264);
   U1365 : MUX2_X1 port map( A => n1215, B => n308, S => n484, Z => n3263);
   U1366 : MUX2_X1 port map( A => n1216, B => n311, S => n483, Z => n3262);
   U1367 : MUX2_X1 port map( A => n1217, B => n314, S => n483, Z => n3261);
   U1368 : MUX2_X1 port map( A => n1218, B => n317, S => n483, Z => n3260);
   U1369 : MUX2_X1 port map( A => n1219, B => n320, S => n483, Z => n3259);
   U1370 : MUX2_X1 port map( A => n1220, B => n323, S => n483, Z => n3258);
   U1371 : MUX2_X1 port map( A => n1221, B => n326, S => n483, Z => n3257);
   U1372 : MUX2_X1 port map( A => n1222, B => n329, S => n483, Z => n3256);
   U1373 : MUX2_X1 port map( A => n1223, B => n332, S => n483, Z => n3255);
   U1374 : MUX2_X1 port map( A => n1224, B => n335, S => n483, Z => n3254);
   U1375 : MUX2_X1 port map( A => n1225, B => n338, S => n483, Z => n3253);
   U1376 : MUX2_X1 port map( A => n1226, B => n341, S => n483, Z => n3252);
   U1377 : MUX2_X1 port map( A => n1227, B => n344, S => n483, Z => n3251);
   U1378 : MUX2_X1 port map( A => n1228, B => n347, S => n482, Z => n3250);
   U1379 : MUX2_X1 port map( A => n1229, B => n350, S => n482, Z => n3249);
   U1380 : MUX2_X1 port map( A => n1230, B => n353, S => n482, Z => n3248);
   U1381 : MUX2_X1 port map( A => n1231, B => n356, S => n482, Z => n3247);
   U1382 : MUX2_X1 port map( A => n1232, B => n359, S => n482, Z => n3246);
   U1383 : MUX2_X1 port map( A => n1233, B => n362, S => n482, Z => n3245);
   U1384 : MUX2_X1 port map( A => n1234, B => n365, S => n482, Z => n3244);
   U1385 : MUX2_X1 port map( A => n1235, B => n368, S => n482, Z => n3243);
   U1386 : MUX2_X1 port map( A => n1236, B => n371, S => n482, Z => n3242);
   U1387 : MUX2_X1 port map( A => n1237, B => n374, S => n482, Z => n3241);
   U1388 : MUX2_X1 port map( A => n1238, B => n377, S => n482, Z => n3240);
   U1389 : MUX2_X1 port map( A => n1239, B => n380, S => n482, Z => n3239);
   U1390 : OAI21_X1 port map( B1 => n851, B2 => n1205, A => n260, ZN => n1208);
   U1391 : MUX2_X1 port map( A => n1240, B => n283, S => n488, Z => n3238);
   U1392 : MUX2_X1 port map( A => n1242, B => n290, S => n488, Z => n3237);
   U1393 : MUX2_X1 port map( A => n1243, B => n293, S => n488, Z => n3236);
   U1394 : MUX2_X1 port map( A => n1244, B => n296, S => n488, Z => n3235);
   U1395 : MUX2_X1 port map( A => n1245, B => n299, S => n488, Z => n3234);
   U1396 : MUX2_X1 port map( A => n1246, B => n302, S => n488, Z => n3233);
   U1397 : MUX2_X1 port map( A => n1247, B => n305, S => n488, Z => n3232);
   U1398 : MUX2_X1 port map( A => n1248, B => n308, S => n488, Z => n3231);
   U1399 : MUX2_X1 port map( A => n1249, B => n311, S => n487, Z => n3230);
   U1400 : MUX2_X1 port map( A => n1250, B => n314, S => n487, Z => n3229);
   U1401 : MUX2_X1 port map( A => n1251, B => n317, S => n487, Z => n3228);
   U1402 : MUX2_X1 port map( A => n1252, B => n320, S => n487, Z => n3227);
   U1403 : MUX2_X1 port map( A => n1253, B => n323, S => n487, Z => n3226);
   U1404 : MUX2_X1 port map( A => n1254, B => n326, S => n487, Z => n3225);
   U1405 : MUX2_X1 port map( A => n1255, B => n329, S => n487, Z => n3224);
   U1406 : MUX2_X1 port map( A => n1256, B => n332, S => n487, Z => n3223);
   U1407 : MUX2_X1 port map( A => n1257, B => n335, S => n487, Z => n3222);
   U1408 : MUX2_X1 port map( A => n1258, B => n338, S => n487, Z => n3221);
   U1409 : MUX2_X1 port map( A => n1259, B => n341, S => n487, Z => n3220);
   U1410 : MUX2_X1 port map( A => n1260, B => n344, S => n487, Z => n3219);
   U1411 : MUX2_X1 port map( A => n1261, B => n347, S => n486, Z => n3218);
   U1412 : MUX2_X1 port map( A => n1262, B => n350, S => n486, Z => n3217);
   U1413 : MUX2_X1 port map( A => n1263, B => n353, S => n486, Z => n3216);
   U1414 : MUX2_X1 port map( A => n1264, B => n356, S => n486, Z => n3215);
   U1415 : MUX2_X1 port map( A => n1265, B => n359, S => n486, Z => n3214);
   U1416 : MUX2_X1 port map( A => n1266, B => n362, S => n486, Z => n3213);
   U1417 : MUX2_X1 port map( A => n1267, B => n365, S => n486, Z => n3212);
   U1418 : MUX2_X1 port map( A => n1268, B => n368, S => n486, Z => n3211);
   U1419 : MUX2_X1 port map( A => n1269, B => n371, S => n486, Z => n3210);
   U1420 : MUX2_X1 port map( A => n1270, B => n374, S => n486, Z => n3209);
   U1421 : MUX2_X1 port map( A => n1271, B => n377, S => n486, Z => n3208);
   U1422 : MUX2_X1 port map( A => n1272, B => n380, S => n486, Z => n3207);
   U1423 : OAI21_X1 port map( B1 => n853, B2 => n1205, A => n262, ZN => n1241);
   U1424 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => n854, A3 => n1134, ZN => 
                           n1205);
   U1425 : INV_X1 port map( A => ADD_WR(2), ZN => n854);
   U1426 : MUX2_X1 port map( A => n4467, B => n283, S => n492, Z => n3206);
   U1427 : MUX2_X1 port map( A => n4466, B => n290, S => n492, Z => n3205);
   U1428 : MUX2_X1 port map( A => n4465, B => n293, S => n492, Z => n3204);
   U1429 : MUX2_X1 port map( A => n4464, B => n296, S => n492, Z => n3203);
   U1430 : MUX2_X1 port map( A => n4463, B => n299, S => n492, Z => n3202);
   U1431 : MUX2_X1 port map( A => n4462, B => n302, S => n492, Z => n3201);
   U1432 : MUX2_X1 port map( A => n4461, B => n305, S => n492, Z => n3200);
   U1433 : MUX2_X1 port map( A => n4460, B => n308, S => n492, Z => n3199);
   U1434 : MUX2_X1 port map( A => n4459, B => n311, S => n491, Z => n3198);
   U1435 : MUX2_X1 port map( A => n4458, B => n314, S => n491, Z => n3197);
   U1436 : MUX2_X1 port map( A => n4457, B => n317, S => n491, Z => n3196);
   U1437 : MUX2_X1 port map( A => n4456, B => n320, S => n491, Z => n3195);
   U1438 : MUX2_X1 port map( A => n4455, B => n323, S => n491, Z => n3194);
   U1439 : MUX2_X1 port map( A => n4454, B => n326, S => n491, Z => n3193);
   U1440 : MUX2_X1 port map( A => n4453, B => n329, S => n491, Z => n3192);
   U1441 : MUX2_X1 port map( A => n4452, B => n332, S => n491, Z => n3191);
   U1442 : MUX2_X1 port map( A => n4451, B => n335, S => n491, Z => n3190);
   U1443 : MUX2_X1 port map( A => n4450, B => n338, S => n491, Z => n3189);
   U1444 : MUX2_X1 port map( A => n4449, B => n341, S => n491, Z => n3188);
   U1445 : MUX2_X1 port map( A => n4448, B => n344, S => n491, Z => n3187);
   U1446 : MUX2_X1 port map( A => n4447, B => n347, S => n490, Z => n3186);
   U1447 : MUX2_X1 port map( A => n4446, B => n350, S => n490, Z => n3185);
   U1448 : MUX2_X1 port map( A => n4445, B => n353, S => n490, Z => n3184);
   U1449 : MUX2_X1 port map( A => n4444, B => n356, S => n490, Z => n3183);
   U1450 : MUX2_X1 port map( A => n4443, B => n359, S => n490, Z => n3182);
   U1451 : MUX2_X1 port map( A => n4442, B => n362, S => n490, Z => n3181);
   U1452 : MUX2_X1 port map( A => n4441, B => n365, S => n490, Z => n3180);
   U1453 : MUX2_X1 port map( A => n4440, B => n368, S => n490, Z => n3179);
   U1454 : MUX2_X1 port map( A => n4439, B => n371, S => n490, Z => n3178);
   U1455 : MUX2_X1 port map( A => n4438, B => n374, S => n490, Z => n3177);
   U1456 : MUX2_X1 port map( A => n4437, B => n377, S => n490, Z => n3176);
   U1457 : MUX2_X1 port map( A => n4436, B => n380, S => n490, Z => n3175);
   U1458 : OAI21_X1 port map( B1 => n815, B2 => n1274, A => n262, ZN => n1273);
   U1459 : NAND2_X1 port map( A1 => n1275, A2 => n1276, ZN => n815);
   U1460 : MUX2_X1 port map( A => n4435, B => n283, S => n496, Z => n3174);
   U1461 : MUX2_X1 port map( A => n4434, B => n290, S => n496, Z => n3173);
   U1462 : MUX2_X1 port map( A => n4433, B => n293, S => n496, Z => n3172);
   U1463 : MUX2_X1 port map( A => n4432, B => n296, S => n496, Z => n3171);
   U1464 : MUX2_X1 port map( A => n4431, B => n299, S => n496, Z => n3170);
   U1465 : MUX2_X1 port map( A => n4430, B => n302, S => n496, Z => n3169);
   U1466 : MUX2_X1 port map( A => n4429, B => n305, S => n496, Z => n3168);
   U1467 : MUX2_X1 port map( A => n4428, B => n308, S => n496, Z => n3167);
   U1468 : MUX2_X1 port map( A => n4427, B => n311, S => n495, Z => n3166);
   U1469 : MUX2_X1 port map( A => n4426, B => n314, S => n495, Z => n3165);
   U1470 : MUX2_X1 port map( A => n4425, B => n317, S => n495, Z => n3164);
   U1471 : MUX2_X1 port map( A => n4424, B => n320, S => n495, Z => n3163);
   U1472 : MUX2_X1 port map( A => n4423, B => n323, S => n495, Z => n3162);
   U1473 : MUX2_X1 port map( A => n4422, B => n326, S => n495, Z => n3161);
   U1474 : MUX2_X1 port map( A => n4421, B => n329, S => n495, Z => n3160);
   U1475 : MUX2_X1 port map( A => n4420, B => n332, S => n495, Z => n3159);
   U1476 : MUX2_X1 port map( A => n4419, B => n335, S => n495, Z => n3158);
   U1477 : MUX2_X1 port map( A => n4418, B => n338, S => n495, Z => n3157);
   U1478 : MUX2_X1 port map( A => n4417, B => n341, S => n495, Z => n3156);
   U1479 : MUX2_X1 port map( A => n4416, B => n344, S => n495, Z => n3155);
   U1480 : MUX2_X1 port map( A => n4415, B => n347, S => n494, Z => n3154);
   U1481 : MUX2_X1 port map( A => n4414, B => n350, S => n494, Z => n3153);
   U1482 : MUX2_X1 port map( A => n4413, B => n353, S => n494, Z => n3152);
   U1483 : MUX2_X1 port map( A => n4412, B => n356, S => n494, Z => n3151);
   U1484 : MUX2_X1 port map( A => n4411, B => n359, S => n494, Z => n3150);
   U1485 : MUX2_X1 port map( A => n4410, B => n362, S => n494, Z => n3149);
   U1486 : MUX2_X1 port map( A => n4409, B => n365, S => n494, Z => n3148);
   U1487 : MUX2_X1 port map( A => n4408, B => n368, S => n494, Z => n3147);
   U1488 : MUX2_X1 port map( A => n4407, B => n371, S => n494, Z => n3146);
   U1489 : MUX2_X1 port map( A => n4406, B => n374, S => n494, Z => n3145);
   U1490 : MUX2_X1 port map( A => n4405, B => n377, S => n494, Z => n3144);
   U1491 : MUX2_X1 port map( A => n4404, B => n380, S => n494, Z => n3143);
   U1492 : OAI21_X1 port map( B1 => n849, B2 => n1274, A => n262, ZN => n1277);
   U1493 : NAND2_X1 port map( A1 => ADD_WR(0), A2 => n1275, ZN => n849);
   U1494 : INV_X1 port map( A => ADD_WR(1), ZN => n1275);
   U1495 : MUX2_X1 port map( A => n1278, B => n283, S => n500, Z => n3142);
   U1496 : MUX2_X1 port map( A => n1280, B => n290, S => n500, Z => n3141);
   U1497 : MUX2_X1 port map( A => n1281, B => n293, S => n500, Z => n3140);
   U1498 : MUX2_X1 port map( A => n1282, B => n296, S => n500, Z => n3139);
   U1499 : MUX2_X1 port map( A => n1283, B => n299, S => n500, Z => n3138);
   U1500 : MUX2_X1 port map( A => n1284, B => n302, S => n500, Z => n3137);
   U1501 : MUX2_X1 port map( A => n1285, B => n305, S => n500, Z => n3136);
   U1502 : MUX2_X1 port map( A => n1286, B => n308, S => n500, Z => n3135);
   U1503 : MUX2_X1 port map( A => n1287, B => n311, S => n499, Z => n3134);
   U1504 : MUX2_X1 port map( A => n1288, B => n314, S => n499, Z => n3133);
   U1505 : MUX2_X1 port map( A => n1289, B => n317, S => n499, Z => n3132);
   U1506 : MUX2_X1 port map( A => n1290, B => n320, S => n499, Z => n3131);
   U1507 : MUX2_X1 port map( A => n1291, B => n323, S => n499, Z => n3130);
   U1508 : MUX2_X1 port map( A => n1292, B => n326, S => n499, Z => n3129);
   U1509 : MUX2_X1 port map( A => n1293, B => n329, S => n499, Z => n3128);
   U1510 : MUX2_X1 port map( A => n1294, B => n332, S => n499, Z => n3127);
   U1511 : MUX2_X1 port map( A => n1295, B => n335, S => n499, Z => n3126);
   U1512 : MUX2_X1 port map( A => n1296, B => n338, S => n499, Z => n3125);
   U1513 : MUX2_X1 port map( A => n1297, B => n341, S => n499, Z => n3124);
   U1514 : MUX2_X1 port map( A => n1298, B => n344, S => n499, Z => n3123);
   U1515 : MUX2_X1 port map( A => n1299, B => n347, S => n498, Z => n3122);
   U1516 : MUX2_X1 port map( A => n1300, B => n350, S => n498, Z => n3121);
   U1517 : MUX2_X1 port map( A => n1301, B => n353, S => n498, Z => n3120);
   U1518 : MUX2_X1 port map( A => n1302, B => n356, S => n498, Z => n3119);
   U1519 : MUX2_X1 port map( A => n1303, B => n359, S => n498, Z => n3118);
   U1520 : MUX2_X1 port map( A => n1304, B => n362, S => n498, Z => n3117);
   U1521 : MUX2_X1 port map( A => n1305, B => n365, S => n498, Z => n3116);
   U1522 : MUX2_X1 port map( A => n1306, B => n368, S => n498, Z => n3115);
   U1523 : MUX2_X1 port map( A => n1307, B => n371, S => n498, Z => n3114);
   U1524 : MUX2_X1 port map( A => n1308, B => n374, S => n498, Z => n3113);
   U1525 : MUX2_X1 port map( A => n1309, B => n377, S => n498, Z => n3112);
   U1526 : MUX2_X1 port map( A => n1310, B => n380, S => n498, Z => n3111);
   U1527 : OAI21_X1 port map( B1 => n851, B2 => n1274, A => n262, ZN => n1279);
   U1528 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => n1276, ZN => n851);
   U1529 : INV_X1 port map( A => ADD_WR(0), ZN => n1276);
   U1530 : MUX2_X1 port map( A => n1311, B => n283, S => n504, Z => n3110);
   U1531 : INV_X1 port map( A => n1313, ZN => n750);
   U1532 : OAI221_X1 port map( B1 => n1313, B2 => n505, C1 => n275, C2 => n1315
                           , A => n1316, ZN => n3109);
   U1533 : OAI21_X1 port map( B1 => n1317, B2 => n1318, A => n510, ZN => n1316)
                           ;
   U1534 : NAND4_X1 port map( A1 => n1320, A2 => n1321, A3 => n1322, A4 => 
                           n1323, ZN => n1318);
   U1535 : AOI221_X1 port map( B1 => n513, B2 => n1029, C1 => n516, C2 => n995,
                           A => n1326, ZN => n1323);
   U1536 : OAI22_X1 port map( A1 => n5075, A2 => n519, B1 => n5107, B2 => n522,
                           ZN => n1326);
   U1537 : AOI221_X1 port map( B1 => n525, B2 => n857, C1 => n528, C2 => n891, 
                           A => n1331, ZN => n1322);
   U1538 : OAI22_X1 port map( A1 => n5363, A2 => n531, B1 => n5331, B2 => n534,
                           ZN => n1331);
   U1539 : AOI221_X1 port map( B1 => n537, B2 => n1311, C1 => n540, C2 => n1278
                           , A => n1336, ZN => n1321);
   U1540 : OAI22_X1 port map( A1 => n4499, A2 => n543, B1 => n4531, B2 => n546,
                           ZN => n1336);
   U1541 : AOI221_X1 port map( B1 => n549, B2 => n1099, C1 => n552, C2 => n1065
                           , A => n1341, ZN => n1320);
   U1542 : OAI22_X1 port map( A1 => n4691, A2 => n555, B1 => n4723, B2 => n558,
                           ZN => n1341);
   U1543 : NAND4_X1 port map( A1 => n1344, A2 => n1345, A3 => n1346, A4 => 
                           n1347, ZN => n1317);
   U1544 : AOI221_X1 port map( B1 => n561, B2 => n5011, C1 => n564, C2 => n5043
                           , A => n1350, ZN => n1347);
   U1545 : OAI22_X1 port map( A1 => n1351, A2 => n567, B1 => n1353, B2 => n570,
                           ZN => n1350);
   U1546 : AOI221_X1 port map( B1 => n573, B2 => n5299, C1 => n576, C2 => n5267
                           , A => n1357, ZN => n1346);
   U1547 : OAI22_X1 port map( A1 => n1358, A2 => n579, B1 => n1360, B2 => n582,
                           ZN => n1357);
   U1548 : AOI221_X1 port map( B1 => n585, B2 => n4563, C1 => n588, C2 => n4595
                           , A => n1364, ZN => n1345);
   U1549 : OAI22_X1 port map( A1 => n1365, A2 => n591, B1 => n1367, B2 => n594,
                           ZN => n1364);
   U1550 : AOI221_X1 port map( B1 => n597, B2 => n4627, C1 => n600, C2 => n4659
                           , A => n1371, ZN => n1344);
   U1551 : OAI22_X1 port map( A1 => n1372, A2 => n603, B1 => n1374, B2 => n606,
                           ZN => n1371);
   U1552 : MUX2_X1 port map( A => n1376, B => n290, S => n504, Z => n3108);
   U1553 : INV_X1 port map( A => n1377, ZN => n753);
   U1554 : OAI221_X1 port map( B1 => n1377, B2 => n505, C1 => n272, C2 => n1378
                           , A => n1379, ZN => n3107);
   U1555 : OAI21_X1 port map( B1 => n1380, B2 => n1381, A => n510, ZN => n1379)
                           ;
   U1556 : NAND4_X1 port map( A1 => n1382, A2 => n1383, A3 => n1384, A4 => 
                           n1385, ZN => n1381);
   U1557 : AOI221_X1 port map( B1 => n513, B2 => n1031, C1 => n516, C2 => n997,
                           A => n1386, ZN => n1385);
   U1558 : OAI22_X1 port map( A1 => n5074, A2 => n519, B1 => n5106, B2 => n522,
                           ZN => n1386);
   U1559 : AOI221_X1 port map( B1 => n525, B2 => n859, C1 => n528, C2 => n893, 
                           A => n1387, ZN => n1384);
   U1560 : OAI22_X1 port map( A1 => n5362, A2 => n531, B1 => n5330, B2 => n534,
                           ZN => n1387);
   U1561 : AOI221_X1 port map( B1 => n537, B2 => n1376, C1 => n540, C2 => n1280
                           , A => n1388, ZN => n1383);
   U1562 : OAI22_X1 port map( A1 => n4498, A2 => n543, B1 => n4530, B2 => n546,
                           ZN => n1388);
   U1563 : AOI221_X1 port map( B1 => n549, B2 => n1101, C1 => n552, C2 => n1067
                           , A => n1389, ZN => n1382);
   U1564 : OAI22_X1 port map( A1 => n4690, A2 => n555, B1 => n4722, B2 => n558,
                           ZN => n1389);
   U1565 : NAND4_X1 port map( A1 => n1390, A2 => n1391, A3 => n1392, A4 => 
                           n1393, ZN => n1380);
   U1566 : AOI221_X1 port map( B1 => n561, B2 => n5010, C1 => n564, C2 => n5042
                           , A => n1394, ZN => n1393);
   U1567 : OAI22_X1 port map( A1 => n1395, A2 => n567, B1 => n1396, B2 => n570,
                           ZN => n1394);
   U1568 : AOI221_X1 port map( B1 => n573, B2 => n5298, C1 => n576, C2 => n5266
                           , A => n1397, ZN => n1392);
   U1569 : OAI22_X1 port map( A1 => n1398, A2 => n579, B1 => n1399, B2 => n582,
                           ZN => n1397);
   U1570 : AOI221_X1 port map( B1 => n585, B2 => n4562, C1 => n588, C2 => n4594
                           , A => n1400, ZN => n1391);
   U1571 : OAI22_X1 port map( A1 => n1401, A2 => n591, B1 => n1402, B2 => n594,
                           ZN => n1400);
   U1572 : AOI221_X1 port map( B1 => n597, B2 => n4626, C1 => n600, C2 => n4658
                           , A => n1403, ZN => n1390);
   U1573 : OAI22_X1 port map( A1 => n1404, A2 => n603, B1 => n1405, B2 => n606,
                           ZN => n1403);
   U1574 : MUX2_X1 port map( A => n1406, B => n293, S => n504, Z => n3106);
   U1575 : INV_X1 port map( A => n1407, ZN => n755);
   U1576 : OAI221_X1 port map( B1 => n1407, B2 => n505, C1 => n272, C2 => n1408
                           , A => n1409, ZN => n3105);
   U1577 : OAI21_X1 port map( B1 => n1410, B2 => n1411, A => n510, ZN => n1409)
                           ;
   U1578 : NAND4_X1 port map( A1 => n1412, A2 => n1413, A3 => n1414, A4 => 
                           n1415, ZN => n1411);
   U1579 : AOI221_X1 port map( B1 => n513, B2 => n1032, C1 => n516, C2 => n998,
                           A => n1416, ZN => n1415);
   U1580 : OAI22_X1 port map( A1 => n5073, A2 => n519, B1 => n5105, B2 => n522,
                           ZN => n1416);
   U1581 : AOI221_X1 port map( B1 => n525, B2 => n860, C1 => n528, C2 => n894, 
                           A => n1417, ZN => n1414);
   U1582 : OAI22_X1 port map( A1 => n5361, A2 => n531, B1 => n5329, B2 => n534,
                           ZN => n1417);
   U1583 : AOI221_X1 port map( B1 => n537, B2 => n1406, C1 => n540, C2 => n1281
                           , A => n1418, ZN => n1413);
   U1584 : OAI22_X1 port map( A1 => n4497, A2 => n543, B1 => n4529, B2 => n546,
                           ZN => n1418);
   U1585 : AOI221_X1 port map( B1 => n549, B2 => n1102, C1 => n552, C2 => n1068
                           , A => n1419, ZN => n1412);
   U1586 : OAI22_X1 port map( A1 => n4689, A2 => n555, B1 => n4721, B2 => n558,
                           ZN => n1419);
   U1587 : NAND4_X1 port map( A1 => n1420, A2 => n1421, A3 => n1422, A4 => 
                           n1423, ZN => n1410);
   U1588 : AOI221_X1 port map( B1 => n561, B2 => n5009, C1 => n564, C2 => n5041
                           , A => n1424, ZN => n1423);
   U1589 : OAI22_X1 port map( A1 => n1425, A2 => n567, B1 => n1426, B2 => n570,
                           ZN => n1424);
   U1590 : AOI221_X1 port map( B1 => n573, B2 => n5297, C1 => n576, C2 => n5265
                           , A => n1427, ZN => n1422);
   U1591 : OAI22_X1 port map( A1 => n1428, A2 => n579, B1 => n1429, B2 => n582,
                           ZN => n1427);
   U1592 : AOI221_X1 port map( B1 => n585, B2 => n4561, C1 => n588, C2 => n4593
                           , A => n1430, ZN => n1421);
   U1593 : OAI22_X1 port map( A1 => n1431, A2 => n591, B1 => n1432, B2 => n594,
                           ZN => n1430);
   U1594 : AOI221_X1 port map( B1 => n597, B2 => n4625, C1 => n600, C2 => n4657
                           , A => n1433, ZN => n1420);
   U1595 : OAI22_X1 port map( A1 => n1434, A2 => n603, B1 => n1435, B2 => n606,
                           ZN => n1433);
   U1596 : MUX2_X1 port map( A => n1436, B => n296, S => n504, Z => n3104);
   U1597 : INV_X1 port map( A => n1437, ZN => n757);
   U1598 : OAI221_X1 port map( B1 => n1437, B2 => n505, C1 => n272, C2 => n1438
                           , A => n1439, ZN => n3103);
   U1599 : OAI21_X1 port map( B1 => n1440, B2 => n1441, A => n510, ZN => n1439)
                           ;
   U1600 : NAND4_X1 port map( A1 => n1442, A2 => n1443, A3 => n1444, A4 => 
                           n1445, ZN => n1441);
   U1601 : AOI221_X1 port map( B1 => n513, B2 => n1033, C1 => n516, C2 => n999,
                           A => n1446, ZN => n1445);
   U1602 : OAI22_X1 port map( A1 => n5072, A2 => n519, B1 => n5104, B2 => n522,
                           ZN => n1446);
   U1603 : AOI221_X1 port map( B1 => n525, B2 => n861, C1 => n528, C2 => n895, 
                           A => n1447, ZN => n1444);
   U1604 : OAI22_X1 port map( A1 => n5360, A2 => n531, B1 => n5328, B2 => n534,
                           ZN => n1447);
   U1605 : AOI221_X1 port map( B1 => n537, B2 => n1436, C1 => n540, C2 => n1282
                           , A => n1448, ZN => n1443);
   U1606 : OAI22_X1 port map( A1 => n4496, A2 => n543, B1 => n4528, B2 => n546,
                           ZN => n1448);
   U1607 : AOI221_X1 port map( B1 => n549, B2 => n1103, C1 => n552, C2 => n1069
                           , A => n1449, ZN => n1442);
   U1608 : OAI22_X1 port map( A1 => n4688, A2 => n555, B1 => n4720, B2 => n558,
                           ZN => n1449);
   U1609 : NAND4_X1 port map( A1 => n1450, A2 => n1451, A3 => n1452, A4 => 
                           n1453, ZN => n1440);
   U1610 : AOI221_X1 port map( B1 => n561, B2 => n5008, C1 => n564, C2 => n5040
                           , A => n1454, ZN => n1453);
   U1611 : OAI22_X1 port map( A1 => n1455, A2 => n567, B1 => n1456, B2 => n570,
                           ZN => n1454);
   U1612 : AOI221_X1 port map( B1 => n573, B2 => n5296, C1 => n576, C2 => n5264
                           , A => n1457, ZN => n1452);
   U1613 : OAI22_X1 port map( A1 => n1458, A2 => n579, B1 => n1459, B2 => n582,
                           ZN => n1457);
   U1614 : AOI221_X1 port map( B1 => n585, B2 => n4560, C1 => n588, C2 => n4592
                           , A => n1460, ZN => n1451);
   U1615 : OAI22_X1 port map( A1 => n1461, A2 => n591, B1 => n1462, B2 => n594,
                           ZN => n1460);
   U1616 : AOI221_X1 port map( B1 => n597, B2 => n4624, C1 => n600, C2 => n4656
                           , A => n1463, ZN => n1450);
   U1617 : OAI22_X1 port map( A1 => n1464, A2 => n603, B1 => n1465, B2 => n606,
                           ZN => n1463);
   U1618 : MUX2_X1 port map( A => n1466, B => n299, S => n504, Z => n3102);
   U1619 : INV_X1 port map( A => n1467, ZN => n759);
   U1620 : OAI221_X1 port map( B1 => n1467, B2 => n505, C1 => n274, C2 => n1468
                           , A => n1469, ZN => n3101);
   U1621 : OAI21_X1 port map( B1 => n1470, B2 => n1471, A => n510, ZN => n1469)
                           ;
   U1622 : NAND4_X1 port map( A1 => n1472, A2 => n1473, A3 => n1474, A4 => 
                           n1475, ZN => n1471);
   U1623 : AOI221_X1 port map( B1 => n513, B2 => n1034, C1 => n516, C2 => n1000
                           , A => n1476, ZN => n1475);
   U1624 : OAI22_X1 port map( A1 => n5071, A2 => n519, B1 => n5103, B2 => n522,
                           ZN => n1476);
   U1625 : AOI221_X1 port map( B1 => n525, B2 => n862, C1 => n528, C2 => n896, 
                           A => n1477, ZN => n1474);
   U1626 : OAI22_X1 port map( A1 => n5359, A2 => n531, B1 => n5327, B2 => n534,
                           ZN => n1477);
   U1627 : AOI221_X1 port map( B1 => n537, B2 => n1466, C1 => n540, C2 => n1283
                           , A => n1478, ZN => n1473);
   U1628 : OAI22_X1 port map( A1 => n4495, A2 => n543, B1 => n4527, B2 => n546,
                           ZN => n1478);
   U1629 : AOI221_X1 port map( B1 => n549, B2 => n1104, C1 => n552, C2 => n1070
                           , A => n1479, ZN => n1472);
   U1630 : OAI22_X1 port map( A1 => n4687, A2 => n555, B1 => n4719, B2 => n558,
                           ZN => n1479);
   U1631 : NAND4_X1 port map( A1 => n1480, A2 => n1481, A3 => n1482, A4 => 
                           n1483, ZN => n1470);
   U1632 : AOI221_X1 port map( B1 => n561, B2 => n5007, C1 => n564, C2 => n5039
                           , A => n1484, ZN => n1483);
   U1633 : OAI22_X1 port map( A1 => n1485, A2 => n567, B1 => n1486, B2 => n570,
                           ZN => n1484);
   U1634 : AOI221_X1 port map( B1 => n573, B2 => n5295, C1 => n576, C2 => n5263
                           , A => n1487, ZN => n1482);
   U1635 : OAI22_X1 port map( A1 => n1488, A2 => n579, B1 => n1489, B2 => n582,
                           ZN => n1487);
   U1636 : AOI221_X1 port map( B1 => n585, B2 => n4559, C1 => n588, C2 => n4591
                           , A => n1490, ZN => n1481);
   U1637 : OAI22_X1 port map( A1 => n1491, A2 => n591, B1 => n1492, B2 => n594,
                           ZN => n1490);
   U1638 : AOI221_X1 port map( B1 => n597, B2 => n4623, C1 => n600, C2 => n4655
                           , A => n1493, ZN => n1480);
   U1639 : OAI22_X1 port map( A1 => n1494, A2 => n603, B1 => n1495, B2 => n606,
                           ZN => n1493);
   U1640 : MUX2_X1 port map( A => n1496, B => n302, S => n504, Z => n3100);
   U1641 : INV_X1 port map( A => n1497, ZN => n761);
   U1642 : OAI221_X1 port map( B1 => n1497, B2 => n505, C1 => n272, C2 => n1498
                           , A => n1499, ZN => n3099);
   U1643 : OAI21_X1 port map( B1 => n1500, B2 => n1501, A => n510, ZN => n1499)
                           ;
   U1644 : NAND4_X1 port map( A1 => n1502, A2 => n1503, A3 => n1504, A4 => 
                           n1505, ZN => n1501);
   U1645 : AOI221_X1 port map( B1 => n513, B2 => n1035, C1 => n516, C2 => n1001
                           , A => n1506, ZN => n1505);
   U1646 : OAI22_X1 port map( A1 => n5070, A2 => n519, B1 => n5102, B2 => n522,
                           ZN => n1506);
   U1647 : AOI221_X1 port map( B1 => n525, B2 => n863, C1 => n528, C2 => n897, 
                           A => n1507, ZN => n1504);
   U1648 : OAI22_X1 port map( A1 => n5358, A2 => n531, B1 => n5326, B2 => n534,
                           ZN => n1507);
   U1649 : AOI221_X1 port map( B1 => n537, B2 => n1496, C1 => n540, C2 => n1284
                           , A => n1508, ZN => n1503);
   U1650 : OAI22_X1 port map( A1 => n4494, A2 => n543, B1 => n4526, B2 => n546,
                           ZN => n1508);
   U1651 : AOI221_X1 port map( B1 => n549, B2 => n1105, C1 => n552, C2 => n1071
                           , A => n1509, ZN => n1502);
   U1652 : OAI22_X1 port map( A1 => n4686, A2 => n555, B1 => n4718, B2 => n558,
                           ZN => n1509);
   U1653 : NAND4_X1 port map( A1 => n1510, A2 => n1511, A3 => n1512, A4 => 
                           n1513, ZN => n1500);
   U1654 : AOI221_X1 port map( B1 => n561, B2 => n5006, C1 => n564, C2 => n5038
                           , A => n1514, ZN => n1513);
   U1655 : OAI22_X1 port map( A1 => n1515, A2 => n567, B1 => n1516, B2 => n570,
                           ZN => n1514);
   U1656 : AOI221_X1 port map( B1 => n573, B2 => n5294, C1 => n576, C2 => n5262
                           , A => n1517, ZN => n1512);
   U1657 : OAI22_X1 port map( A1 => n1518, A2 => n579, B1 => n1519, B2 => n582,
                           ZN => n1517);
   U1658 : AOI221_X1 port map( B1 => n585, B2 => n4558, C1 => n588, C2 => n4590
                           , A => n1520, ZN => n1511);
   U1659 : OAI22_X1 port map( A1 => n1521, A2 => n591, B1 => n1522, B2 => n594,
                           ZN => n1520);
   U1660 : AOI221_X1 port map( B1 => n597, B2 => n4622, C1 => n600, C2 => n4654
                           , A => n1523, ZN => n1510);
   U1661 : OAI22_X1 port map( A1 => n1524, A2 => n603, B1 => n1525, B2 => n606,
                           ZN => n1523);
   U1662 : MUX2_X1 port map( A => n1526, B => n305, S => n504, Z => n3098);
   U1663 : INV_X1 port map( A => n1527, ZN => n763);
   U1664 : OAI221_X1 port map( B1 => n1527, B2 => n505, C1 => n272, C2 => n1528
                           , A => n1529, ZN => n3097);
   U1665 : OAI21_X1 port map( B1 => n1530, B2 => n1531, A => n510, ZN => n1529)
                           ;
   U1666 : NAND4_X1 port map( A1 => n1532, A2 => n1533, A3 => n1534, A4 => 
                           n1535, ZN => n1531);
   U1667 : AOI221_X1 port map( B1 => n513, B2 => n1036, C1 => n516, C2 => n1002
                           , A => n1536, ZN => n1535);
   U1668 : OAI22_X1 port map( A1 => n5069, A2 => n519, B1 => n5101, B2 => n522,
                           ZN => n1536);
   U1669 : AOI221_X1 port map( B1 => n525, B2 => n864, C1 => n528, C2 => n898, 
                           A => n1537, ZN => n1534);
   U1670 : OAI22_X1 port map( A1 => n5357, A2 => n531, B1 => n5325, B2 => n534,
                           ZN => n1537);
   U1671 : AOI221_X1 port map( B1 => n537, B2 => n1526, C1 => n540, C2 => n1285
                           , A => n1538, ZN => n1533);
   U1672 : OAI22_X1 port map( A1 => n4493, A2 => n543, B1 => n4525, B2 => n546,
                           ZN => n1538);
   U1673 : AOI221_X1 port map( B1 => n549, B2 => n1106, C1 => n552, C2 => n1072
                           , A => n1539, ZN => n1532);
   U1674 : OAI22_X1 port map( A1 => n4685, A2 => n555, B1 => n4717, B2 => n558,
                           ZN => n1539);
   U1675 : NAND4_X1 port map( A1 => n1540, A2 => n1541, A3 => n1542, A4 => 
                           n1543, ZN => n1530);
   U1676 : AOI221_X1 port map( B1 => n561, B2 => n5005, C1 => n564, C2 => n5037
                           , A => n1544, ZN => n1543);
   U1677 : OAI22_X1 port map( A1 => n1545, A2 => n567, B1 => n1546, B2 => n570,
                           ZN => n1544);
   U1678 : AOI221_X1 port map( B1 => n573, B2 => n5293, C1 => n576, C2 => n5261
                           , A => n1547, ZN => n1542);
   U1679 : OAI22_X1 port map( A1 => n1548, A2 => n579, B1 => n1549, B2 => n582,
                           ZN => n1547);
   U1680 : AOI221_X1 port map( B1 => n585, B2 => n4557, C1 => n588, C2 => n4589
                           , A => n1550, ZN => n1541);
   U1681 : OAI22_X1 port map( A1 => n1551, A2 => n591, B1 => n1552, B2 => n594,
                           ZN => n1550);
   U1682 : AOI221_X1 port map( B1 => n597, B2 => n4621, C1 => n600, C2 => n4653
                           , A => n1553, ZN => n1540);
   U1683 : OAI22_X1 port map( A1 => n1554, A2 => n603, B1 => n1555, B2 => n606,
                           ZN => n1553);
   U1684 : MUX2_X1 port map( A => n1556, B => n308, S => n504, Z => n3096);
   U1685 : INV_X1 port map( A => n1557, ZN => n765);
   U1686 : OAI221_X1 port map( B1 => n1557, B2 => n505, C1 => n272, C2 => n1558
                           , A => n1559, ZN => n3095);
   U1687 : OAI21_X1 port map( B1 => n1560, B2 => n1561, A => n510, ZN => n1559)
                           ;
   U1688 : NAND4_X1 port map( A1 => n1562, A2 => n1563, A3 => n1564, A4 => 
                           n1565, ZN => n1561);
   U1689 : AOI221_X1 port map( B1 => n513, B2 => n1037, C1 => n516, C2 => n1003
                           , A => n1566, ZN => n1565);
   U1690 : OAI22_X1 port map( A1 => n5068, A2 => n519, B1 => n5100, B2 => n522,
                           ZN => n1566);
   U1691 : AOI221_X1 port map( B1 => n525, B2 => n865, C1 => n528, C2 => n899, 
                           A => n1567, ZN => n1564);
   U1692 : OAI22_X1 port map( A1 => n5356, A2 => n531, B1 => n5324, B2 => n534,
                           ZN => n1567);
   U1693 : AOI221_X1 port map( B1 => n537, B2 => n1556, C1 => n540, C2 => n1286
                           , A => n1568, ZN => n1563);
   U1694 : OAI22_X1 port map( A1 => n4492, A2 => n543, B1 => n4524, B2 => n546,
                           ZN => n1568);
   U1695 : AOI221_X1 port map( B1 => n549, B2 => n1107, C1 => n552, C2 => n1073
                           , A => n1569, ZN => n1562);
   U1696 : OAI22_X1 port map( A1 => n4684, A2 => n555, B1 => n4716, B2 => n558,
                           ZN => n1569);
   U1697 : NAND4_X1 port map( A1 => n1570, A2 => n1571, A3 => n1572, A4 => 
                           n1573, ZN => n1560);
   U1698 : AOI221_X1 port map( B1 => n561, B2 => n5004, C1 => n564, C2 => n5036
                           , A => n1574, ZN => n1573);
   U1699 : OAI22_X1 port map( A1 => n1575, A2 => n567, B1 => n1576, B2 => n570,
                           ZN => n1574);
   U1700 : AOI221_X1 port map( B1 => n573, B2 => n5292, C1 => n576, C2 => n5260
                           , A => n1577, ZN => n1572);
   U1701 : OAI22_X1 port map( A1 => n1578, A2 => n579, B1 => n1579, B2 => n582,
                           ZN => n1577);
   U1702 : AOI221_X1 port map( B1 => n585, B2 => n4556, C1 => n588, C2 => n4588
                           , A => n1580, ZN => n1571);
   U1703 : OAI22_X1 port map( A1 => n1581, A2 => n591, B1 => n1582, B2 => n594,
                           ZN => n1580);
   U1704 : AOI221_X1 port map( B1 => n597, B2 => n4620, C1 => n600, C2 => n4652
                           , A => n1583, ZN => n1570);
   U1705 : OAI22_X1 port map( A1 => n1584, A2 => n603, B1 => n1585, B2 => n606,
                           ZN => n1583);
   U1706 : MUX2_X1 port map( A => n1586, B => n311, S => n503, Z => n3094);
   U1707 : INV_X1 port map( A => n1587, ZN => n767);
   U1708 : OAI221_X1 port map( B1 => n1587, B2 => n505, C1 => n273, C2 => n1588
                           , A => n1589, ZN => n3093);
   U1709 : OAI21_X1 port map( B1 => n1590, B2 => n1591, A => n509, ZN => n1589)
                           ;
   U1710 : NAND4_X1 port map( A1 => n1592, A2 => n1593, A3 => n1594, A4 => 
                           n1595, ZN => n1591);
   U1711 : AOI221_X1 port map( B1 => n512, B2 => n1038, C1 => n515, C2 => n1004
                           , A => n1596, ZN => n1595);
   U1712 : OAI22_X1 port map( A1 => n5067, A2 => n518, B1 => n5099, B2 => n521,
                           ZN => n1596);
   U1713 : AOI221_X1 port map( B1 => n524, B2 => n866, C1 => n527, C2 => n900, 
                           A => n1597, ZN => n1594);
   U1714 : OAI22_X1 port map( A1 => n5355, A2 => n530, B1 => n5323, B2 => n533,
                           ZN => n1597);
   U1715 : AOI221_X1 port map( B1 => n536, B2 => n1586, C1 => n539, C2 => n1287
                           , A => n1598, ZN => n1593);
   U1716 : OAI22_X1 port map( A1 => n4491, A2 => n542, B1 => n4523, B2 => n545,
                           ZN => n1598);
   U1717 : AOI221_X1 port map( B1 => n548, B2 => n1108, C1 => n551, C2 => n1074
                           , A => n1599, ZN => n1592);
   U1718 : OAI22_X1 port map( A1 => n4683, A2 => n554, B1 => n4715, B2 => n557,
                           ZN => n1599);
   U1719 : NAND4_X1 port map( A1 => n1600, A2 => n1601, A3 => n1602, A4 => 
                           n1603, ZN => n1590);
   U1720 : AOI221_X1 port map( B1 => n560, B2 => n5003, C1 => n563, C2 => n5035
                           , A => n1604, ZN => n1603);
   U1721 : OAI22_X1 port map( A1 => n1605, A2 => n566, B1 => n1606, B2 => n569,
                           ZN => n1604);
   U1722 : AOI221_X1 port map( B1 => n572, B2 => n5291, C1 => n575, C2 => n5259
                           , A => n1607, ZN => n1602);
   U1723 : OAI22_X1 port map( A1 => n1608, A2 => n578, B1 => n1609, B2 => n581,
                           ZN => n1607);
   U1724 : AOI221_X1 port map( B1 => n584, B2 => n4555, C1 => n587, C2 => n4587
                           , A => n1610, ZN => n1601);
   U1725 : OAI22_X1 port map( A1 => n1611, A2 => n590, B1 => n1612, B2 => n593,
                           ZN => n1610);
   U1726 : AOI221_X1 port map( B1 => n596, B2 => n4619, C1 => n599, C2 => n4651
                           , A => n1613, ZN => n1600);
   U1727 : OAI22_X1 port map( A1 => n1614, A2 => n602, B1 => n1615, B2 => n605,
                           ZN => n1613);
   U1728 : MUX2_X1 port map( A => n1616, B => n314, S => n503, Z => n3092);
   U1729 : INV_X1 port map( A => n1617, ZN => n769);
   U1730 : OAI221_X1 port map( B1 => n1617, B2 => n505, C1 => n272, C2 => n1618
                           , A => n1619, ZN => n3091);
   U1731 : OAI21_X1 port map( B1 => n1620, B2 => n1621, A => n509, ZN => n1619)
                           ;
   U1732 : NAND4_X1 port map( A1 => n1622, A2 => n1623, A3 => n1624, A4 => 
                           n1625, ZN => n1621);
   U1733 : AOI221_X1 port map( B1 => n512, B2 => n1039, C1 => n515, C2 => n1005
                           , A => n1626, ZN => n1625);
   U1734 : OAI22_X1 port map( A1 => n5066, A2 => n518, B1 => n5098, B2 => n521,
                           ZN => n1626);
   U1735 : AOI221_X1 port map( B1 => n524, B2 => n867, C1 => n527, C2 => n901, 
                           A => n1627, ZN => n1624);
   U1736 : OAI22_X1 port map( A1 => n5354, A2 => n530, B1 => n5322, B2 => n533,
                           ZN => n1627);
   U1737 : AOI221_X1 port map( B1 => n536, B2 => n1616, C1 => n539, C2 => n1288
                           , A => n1628, ZN => n1623);
   U1738 : OAI22_X1 port map( A1 => n4490, A2 => n542, B1 => n4522, B2 => n545,
                           ZN => n1628);
   U1739 : AOI221_X1 port map( B1 => n548, B2 => n1109, C1 => n551, C2 => n1075
                           , A => n1629, ZN => n1622);
   U1740 : OAI22_X1 port map( A1 => n4682, A2 => n554, B1 => n4714, B2 => n557,
                           ZN => n1629);
   U1741 : NAND4_X1 port map( A1 => n1630, A2 => n1631, A3 => n1632, A4 => 
                           n1633, ZN => n1620);
   U1742 : AOI221_X1 port map( B1 => n560, B2 => n5002, C1 => n563, C2 => n5034
                           , A => n1634, ZN => n1633);
   U1743 : OAI22_X1 port map( A1 => n1635, A2 => n566, B1 => n1636, B2 => n569,
                           ZN => n1634);
   U1744 : AOI221_X1 port map( B1 => n572, B2 => n5290, C1 => n575, C2 => n5258
                           , A => n1637, ZN => n1632);
   U1745 : OAI22_X1 port map( A1 => n1638, A2 => n578, B1 => n1639, B2 => n581,
                           ZN => n1637);
   U1746 : AOI221_X1 port map( B1 => n584, B2 => n4554, C1 => n587, C2 => n4586
                           , A => n1640, ZN => n1631);
   U1747 : OAI22_X1 port map( A1 => n1641, A2 => n590, B1 => n1642, B2 => n593,
                           ZN => n1640);
   U1748 : AOI221_X1 port map( B1 => n596, B2 => n4618, C1 => n599, C2 => n4650
                           , A => n1643, ZN => n1630);
   U1749 : OAI22_X1 port map( A1 => n1644, A2 => n602, B1 => n1645, B2 => n605,
                           ZN => n1643);
   U1750 : MUX2_X1 port map( A => n1646, B => n317, S => n503, Z => n3090);
   U1751 : INV_X1 port map( A => n1647, ZN => n771);
   U1752 : OAI221_X1 port map( B1 => n1647, B2 => n505, C1 => n271, C2 => n1648
                           , A => n1649, ZN => n3089);
   U1753 : OAI21_X1 port map( B1 => n1650, B2 => n1651, A => n509, ZN => n1649)
                           ;
   U1754 : NAND4_X1 port map( A1 => n1652, A2 => n1653, A3 => n1654, A4 => 
                           n1655, ZN => n1651);
   U1755 : AOI221_X1 port map( B1 => n512, B2 => n1040, C1 => n515, C2 => n1006
                           , A => n1656, ZN => n1655);
   U1756 : OAI22_X1 port map( A1 => n5065, A2 => n518, B1 => n5097, B2 => n521,
                           ZN => n1656);
   U1757 : AOI221_X1 port map( B1 => n524, B2 => n868, C1 => n527, C2 => n902, 
                           A => n1657, ZN => n1654);
   U1758 : OAI22_X1 port map( A1 => n5353, A2 => n530, B1 => n5321, B2 => n533,
                           ZN => n1657);
   U1759 : AOI221_X1 port map( B1 => n536, B2 => n1646, C1 => n539, C2 => n1289
                           , A => n1658, ZN => n1653);
   U1760 : OAI22_X1 port map( A1 => n4489, A2 => n542, B1 => n4521, B2 => n545,
                           ZN => n1658);
   U1761 : AOI221_X1 port map( B1 => n548, B2 => n1110, C1 => n551, C2 => n1076
                           , A => n1659, ZN => n1652);
   U1762 : OAI22_X1 port map( A1 => n4681, A2 => n554, B1 => n4713, B2 => n557,
                           ZN => n1659);
   U1763 : NAND4_X1 port map( A1 => n1660, A2 => n1661, A3 => n1662, A4 => 
                           n1663, ZN => n1650);
   U1764 : AOI221_X1 port map( B1 => n560, B2 => n5001, C1 => n563, C2 => n5033
                           , A => n1664, ZN => n1663);
   U1765 : OAI22_X1 port map( A1 => n1665, A2 => n566, B1 => n1666, B2 => n569,
                           ZN => n1664);
   U1766 : AOI221_X1 port map( B1 => n572, B2 => n5289, C1 => n575, C2 => n5257
                           , A => n1667, ZN => n1662);
   U1767 : OAI22_X1 port map( A1 => n1668, A2 => n578, B1 => n1669, B2 => n581,
                           ZN => n1667);
   U1768 : AOI221_X1 port map( B1 => n584, B2 => n4553, C1 => n587, C2 => n4585
                           , A => n1670, ZN => n1661);
   U1769 : OAI22_X1 port map( A1 => n1671, A2 => n590, B1 => n1672, B2 => n593,
                           ZN => n1670);
   U1770 : AOI221_X1 port map( B1 => n596, B2 => n4617, C1 => n599, C2 => n4649
                           , A => n1673, ZN => n1660);
   U1771 : OAI22_X1 port map( A1 => n1674, A2 => n602, B1 => n1675, B2 => n605,
                           ZN => n1673);
   U1772 : MUX2_X1 port map( A => n1676, B => n320, S => n503, Z => n3088);
   U1773 : INV_X1 port map( A => n1677, ZN => n773);
   U1774 : OAI221_X1 port map( B1 => n1677, B2 => n505, C1 => n271, C2 => n1678
                           , A => n1679, ZN => n3087);
   U1775 : OAI21_X1 port map( B1 => n1680, B2 => n1681, A => n509, ZN => n1679)
                           ;
   U1776 : NAND4_X1 port map( A1 => n1682, A2 => n1683, A3 => n1684, A4 => 
                           n1685, ZN => n1681);
   U1777 : AOI221_X1 port map( B1 => n512, B2 => n1041, C1 => n515, C2 => n1007
                           , A => n1686, ZN => n1685);
   U1778 : OAI22_X1 port map( A1 => n5064, A2 => n518, B1 => n5096, B2 => n521,
                           ZN => n1686);
   U1779 : AOI221_X1 port map( B1 => n524, B2 => n869, C1 => n527, C2 => n903, 
                           A => n1687, ZN => n1684);
   U1780 : OAI22_X1 port map( A1 => n5352, A2 => n530, B1 => n5320, B2 => n533,
                           ZN => n1687);
   U1781 : AOI221_X1 port map( B1 => n536, B2 => n1676, C1 => n539, C2 => n1290
                           , A => n1688, ZN => n1683);
   U1782 : OAI22_X1 port map( A1 => n4488, A2 => n542, B1 => n4520, B2 => n545,
                           ZN => n1688);
   U1783 : AOI221_X1 port map( B1 => n548, B2 => n1111, C1 => n551, C2 => n1077
                           , A => n1689, ZN => n1682);
   U1784 : OAI22_X1 port map( A1 => n4680, A2 => n554, B1 => n4712, B2 => n557,
                           ZN => n1689);
   U1785 : NAND4_X1 port map( A1 => n1690, A2 => n1691, A3 => n1692, A4 => 
                           n1693, ZN => n1680);
   U1786 : AOI221_X1 port map( B1 => n560, B2 => n5000, C1 => n563, C2 => n5032
                           , A => n1694, ZN => n1693);
   U1787 : OAI22_X1 port map( A1 => n1695, A2 => n566, B1 => n1696, B2 => n569,
                           ZN => n1694);
   U1788 : AOI221_X1 port map( B1 => n572, B2 => n5288, C1 => n575, C2 => n5256
                           , A => n1697, ZN => n1692);
   U1789 : OAI22_X1 port map( A1 => n1698, A2 => n578, B1 => n1699, B2 => n581,
                           ZN => n1697);
   U1790 : AOI221_X1 port map( B1 => n584, B2 => n4552, C1 => n587, C2 => n4584
                           , A => n1700, ZN => n1691);
   U1791 : OAI22_X1 port map( A1 => n1701, A2 => n590, B1 => n1702, B2 => n593,
                           ZN => n1700);
   U1792 : AOI221_X1 port map( B1 => n596, B2 => n4616, C1 => n599, C2 => n4648
                           , A => n1703, ZN => n1690);
   U1793 : OAI22_X1 port map( A1 => n1704, A2 => n602, B1 => n1705, B2 => n605,
                           ZN => n1703);
   U1794 : MUX2_X1 port map( A => n1706, B => n323, S => n503, Z => n3086);
   U1795 : INV_X1 port map( A => n1707, ZN => n775);
   U1796 : OAI221_X1 port map( B1 => n1707, B2 => n506, C1 => n274, C2 => n1708
                           , A => n1709, ZN => n3085);
   U1797 : OAI21_X1 port map( B1 => n1710, B2 => n1711, A => n509, ZN => n1709)
                           ;
   U1798 : NAND4_X1 port map( A1 => n1712, A2 => n1713, A3 => n1714, A4 => 
                           n1715, ZN => n1711);
   U1799 : AOI221_X1 port map( B1 => n512, B2 => n1042, C1 => n515, C2 => n1008
                           , A => n1716, ZN => n1715);
   U1800 : OAI22_X1 port map( A1 => n5063, A2 => n518, B1 => n5095, B2 => n521,
                           ZN => n1716);
   U1801 : AOI221_X1 port map( B1 => n524, B2 => n870, C1 => n527, C2 => n904, 
                           A => n1717, ZN => n1714);
   U1802 : OAI22_X1 port map( A1 => n5351, A2 => n530, B1 => n5319, B2 => n533,
                           ZN => n1717);
   U1803 : AOI221_X1 port map( B1 => n536, B2 => n1706, C1 => n539, C2 => n1291
                           , A => n1718, ZN => n1713);
   U1804 : OAI22_X1 port map( A1 => n4487, A2 => n542, B1 => n4519, B2 => n545,
                           ZN => n1718);
   U1805 : AOI221_X1 port map( B1 => n548, B2 => n1112, C1 => n551, C2 => n1078
                           , A => n1719, ZN => n1712);
   U1806 : OAI22_X1 port map( A1 => n4679, A2 => n554, B1 => n4711, B2 => n557,
                           ZN => n1719);
   U1807 : NAND4_X1 port map( A1 => n1720, A2 => n1721, A3 => n1722, A4 => 
                           n1723, ZN => n1710);
   U1808 : AOI221_X1 port map( B1 => n560, B2 => n4999, C1 => n563, C2 => n5031
                           , A => n1724, ZN => n1723);
   U1809 : OAI22_X1 port map( A1 => n1725, A2 => n566, B1 => n1726, B2 => n569,
                           ZN => n1724);
   U1810 : AOI221_X1 port map( B1 => n572, B2 => n5287, C1 => n575, C2 => n5255
                           , A => n1727, ZN => n1722);
   U1811 : OAI22_X1 port map( A1 => n1728, A2 => n578, B1 => n1729, B2 => n581,
                           ZN => n1727);
   U1812 : AOI221_X1 port map( B1 => n584, B2 => n4551, C1 => n587, C2 => n4583
                           , A => n1730, ZN => n1721);
   U1813 : OAI22_X1 port map( A1 => n1731, A2 => n590, B1 => n1732, B2 => n593,
                           ZN => n1730);
   U1814 : AOI221_X1 port map( B1 => n596, B2 => n4615, C1 => n599, C2 => n4647
                           , A => n1733, ZN => n1720);
   U1815 : OAI22_X1 port map( A1 => n1734, A2 => n602, B1 => n1735, B2 => n605,
                           ZN => n1733);
   U1816 : MUX2_X1 port map( A => n1736, B => n326, S => n503, Z => n3084);
   U1817 : INV_X1 port map( A => n1737, ZN => n777);
   U1818 : OAI221_X1 port map( B1 => n1737, B2 => n506, C1 => n271, C2 => n1738
                           , A => n1739, ZN => n3083);
   U1819 : OAI21_X1 port map( B1 => n1740, B2 => n1741, A => n509, ZN => n1739)
                           ;
   U1820 : NAND4_X1 port map( A1 => n1742, A2 => n1743, A3 => n1744, A4 => 
                           n1745, ZN => n1741);
   U1821 : AOI221_X1 port map( B1 => n512, B2 => n1043, C1 => n515, C2 => n1009
                           , A => n1746, ZN => n1745);
   U1822 : OAI22_X1 port map( A1 => n5062, A2 => n518, B1 => n5094, B2 => n521,
                           ZN => n1746);
   U1823 : AOI221_X1 port map( B1 => n524, B2 => n871, C1 => n527, C2 => n905, 
                           A => n1747, ZN => n1744);
   U1824 : OAI22_X1 port map( A1 => n5350, A2 => n530, B1 => n5318, B2 => n533,
                           ZN => n1747);
   U1825 : AOI221_X1 port map( B1 => n536, B2 => n1736, C1 => n539, C2 => n1292
                           , A => n1748, ZN => n1743);
   U1826 : OAI22_X1 port map( A1 => n4486, A2 => n542, B1 => n4518, B2 => n545,
                           ZN => n1748);
   U1827 : AOI221_X1 port map( B1 => n548, B2 => n1113, C1 => n551, C2 => n1079
                           , A => n1749, ZN => n1742);
   U1828 : OAI22_X1 port map( A1 => n4678, A2 => n554, B1 => n4710, B2 => n557,
                           ZN => n1749);
   U1829 : NAND4_X1 port map( A1 => n1750, A2 => n1751, A3 => n1752, A4 => 
                           n1753, ZN => n1740);
   U1830 : AOI221_X1 port map( B1 => n560, B2 => n4998, C1 => n563, C2 => n5030
                           , A => n1754, ZN => n1753);
   U1831 : OAI22_X1 port map( A1 => n1755, A2 => n566, B1 => n1756, B2 => n569,
                           ZN => n1754);
   U1832 : AOI221_X1 port map( B1 => n572, B2 => n5286, C1 => n575, C2 => n5254
                           , A => n1757, ZN => n1752);
   U1833 : OAI22_X1 port map( A1 => n1758, A2 => n578, B1 => n1759, B2 => n581,
                           ZN => n1757);
   U1834 : AOI221_X1 port map( B1 => n584, B2 => n4550, C1 => n587, C2 => n4582
                           , A => n1760, ZN => n1751);
   U1835 : OAI22_X1 port map( A1 => n1761, A2 => n590, B1 => n1762, B2 => n593,
                           ZN => n1760);
   U1836 : AOI221_X1 port map( B1 => n596, B2 => n4614, C1 => n599, C2 => n4646
                           , A => n1763, ZN => n1750);
   U1837 : OAI22_X1 port map( A1 => n1764, A2 => n602, B1 => n1765, B2 => n605,
                           ZN => n1763);
   U1838 : MUX2_X1 port map( A => n1766, B => n329, S => n503, Z => n3082);
   U1839 : INV_X1 port map( A => n1767, ZN => n779);
   U1840 : OAI221_X1 port map( B1 => n1767, B2 => n506, C1 => n271, C2 => n1768
                           , A => n1769, ZN => n3081);
   U1841 : OAI21_X1 port map( B1 => n1770, B2 => n1771, A => n509, ZN => n1769)
                           ;
   U1842 : NAND4_X1 port map( A1 => n1772, A2 => n1773, A3 => n1774, A4 => 
                           n1775, ZN => n1771);
   U1843 : AOI221_X1 port map( B1 => n512, B2 => n1044, C1 => n515, C2 => n1010
                           , A => n1776, ZN => n1775);
   U1844 : OAI22_X1 port map( A1 => n5061, A2 => n518, B1 => n5093, B2 => n521,
                           ZN => n1776);
   U1845 : AOI221_X1 port map( B1 => n524, B2 => n872, C1 => n527, C2 => n906, 
                           A => n1777, ZN => n1774);
   U1846 : OAI22_X1 port map( A1 => n5349, A2 => n530, B1 => n5317, B2 => n533,
                           ZN => n1777);
   U1847 : AOI221_X1 port map( B1 => n536, B2 => n1766, C1 => n539, C2 => n1293
                           , A => n1778, ZN => n1773);
   U1848 : OAI22_X1 port map( A1 => n4485, A2 => n542, B1 => n4517, B2 => n545,
                           ZN => n1778);
   U1849 : AOI221_X1 port map( B1 => n548, B2 => n1114, C1 => n551, C2 => n1080
                           , A => n1779, ZN => n1772);
   U1850 : OAI22_X1 port map( A1 => n4677, A2 => n554, B1 => n4709, B2 => n557,
                           ZN => n1779);
   U1851 : NAND4_X1 port map( A1 => n1780, A2 => n1781, A3 => n1782, A4 => 
                           n1783, ZN => n1770);
   U1852 : AOI221_X1 port map( B1 => n560, B2 => n4997, C1 => n563, C2 => n5029
                           , A => n1784, ZN => n1783);
   U1853 : OAI22_X1 port map( A1 => n1785, A2 => n566, B1 => n1786, B2 => n569,
                           ZN => n1784);
   U1854 : AOI221_X1 port map( B1 => n572, B2 => n5285, C1 => n575, C2 => n5253
                           , A => n1787, ZN => n1782);
   U1855 : OAI22_X1 port map( A1 => n1788, A2 => n578, B1 => n1789, B2 => n581,
                           ZN => n1787);
   U1856 : AOI221_X1 port map( B1 => n584, B2 => n4549, C1 => n587, C2 => n4581
                           , A => n1790, ZN => n1781);
   U1857 : OAI22_X1 port map( A1 => n1791, A2 => n590, B1 => n1792, B2 => n593,
                           ZN => n1790);
   U1858 : AOI221_X1 port map( B1 => n596, B2 => n4613, C1 => n599, C2 => n4645
                           , A => n1793, ZN => n1780);
   U1859 : OAI22_X1 port map( A1 => n1794, A2 => n602, B1 => n1795, B2 => n605,
                           ZN => n1793);
   U1860 : MUX2_X1 port map( A => n1796, B => n332, S => n503, Z => n3080);
   U1861 : INV_X1 port map( A => n1797, ZN => n781);
   U1862 : OAI221_X1 port map( B1 => n1797, B2 => n506, C1 => n271, C2 => n1798
                           , A => n1799, ZN => n3079);
   U1863 : OAI21_X1 port map( B1 => n1800, B2 => n1801, A => n509, ZN => n1799)
                           ;
   U1864 : NAND4_X1 port map( A1 => n1802, A2 => n1803, A3 => n1804, A4 => 
                           n1805, ZN => n1801);
   U1865 : AOI221_X1 port map( B1 => n512, B2 => n1045, C1 => n515, C2 => n1011
                           , A => n1806, ZN => n1805);
   U1866 : OAI22_X1 port map( A1 => n5060, A2 => n518, B1 => n5092, B2 => n521,
                           ZN => n1806);
   U1867 : AOI221_X1 port map( B1 => n524, B2 => n873, C1 => n527, C2 => n907, 
                           A => n1807, ZN => n1804);
   U1868 : OAI22_X1 port map( A1 => n5348, A2 => n530, B1 => n5316, B2 => n533,
                           ZN => n1807);
   U1869 : AOI221_X1 port map( B1 => n536, B2 => n1796, C1 => n539, C2 => n1294
                           , A => n1808, ZN => n1803);
   U1870 : OAI22_X1 port map( A1 => n4484, A2 => n542, B1 => n4516, B2 => n545,
                           ZN => n1808);
   U1871 : AOI221_X1 port map( B1 => n548, B2 => n1115, C1 => n551, C2 => n1081
                           , A => n1809, ZN => n1802);
   U1872 : OAI22_X1 port map( A1 => n4676, A2 => n554, B1 => n4708, B2 => n557,
                           ZN => n1809);
   U1873 : NAND4_X1 port map( A1 => n1810, A2 => n1811, A3 => n1812, A4 => 
                           n1813, ZN => n1800);
   U1874 : AOI221_X1 port map( B1 => n560, B2 => n4996, C1 => n563, C2 => n5028
                           , A => n1814, ZN => n1813);
   U1875 : OAI22_X1 port map( A1 => n1815, A2 => n566, B1 => n1816, B2 => n569,
                           ZN => n1814);
   U1876 : AOI221_X1 port map( B1 => n572, B2 => n5284, C1 => n575, C2 => n5252
                           , A => n1817, ZN => n1812);
   U1877 : OAI22_X1 port map( A1 => n1818, A2 => n578, B1 => n1819, B2 => n581,
                           ZN => n1817);
   U1878 : AOI221_X1 port map( B1 => n584, B2 => n4548, C1 => n587, C2 => n4580
                           , A => n1820, ZN => n1811);
   U1879 : OAI22_X1 port map( A1 => n1821, A2 => n590, B1 => n1822, B2 => n593,
                           ZN => n1820);
   U1880 : AOI221_X1 port map( B1 => n596, B2 => n4612, C1 => n599, C2 => n4644
                           , A => n1823, ZN => n1810);
   U1881 : OAI22_X1 port map( A1 => n1824, A2 => n602, B1 => n1825, B2 => n605,
                           ZN => n1823);
   U1882 : MUX2_X1 port map( A => n1826, B => n335, S => n503, Z => n3078);
   U1883 : INV_X1 port map( A => n1827, ZN => n783);
   U1884 : OAI221_X1 port map( B1 => n1827, B2 => n506, C1 => n275, C2 => n1828
                           , A => n1829, ZN => n3077);
   U1885 : OAI21_X1 port map( B1 => n1830, B2 => n1831, A => n509, ZN => n1829)
                           ;
   U1886 : NAND4_X1 port map( A1 => n1832, A2 => n1833, A3 => n1834, A4 => 
                           n1835, ZN => n1831);
   U1887 : AOI221_X1 port map( B1 => n512, B2 => n1046, C1 => n515, C2 => n1012
                           , A => n1836, ZN => n1835);
   U1888 : OAI22_X1 port map( A1 => n5059, A2 => n518, B1 => n5091, B2 => n521,
                           ZN => n1836);
   U1889 : AOI221_X1 port map( B1 => n524, B2 => n874, C1 => n527, C2 => n908, 
                           A => n1837, ZN => n1834);
   U1890 : OAI22_X1 port map( A1 => n5347, A2 => n530, B1 => n5315, B2 => n533,
                           ZN => n1837);
   U1891 : AOI221_X1 port map( B1 => n536, B2 => n1826, C1 => n539, C2 => n1295
                           , A => n1838, ZN => n1833);
   U1892 : OAI22_X1 port map( A1 => n4483, A2 => n542, B1 => n4515, B2 => n545,
                           ZN => n1838);
   U1893 : AOI221_X1 port map( B1 => n548, B2 => n1116, C1 => n551, C2 => n1082
                           , A => n1839, ZN => n1832);
   U1894 : OAI22_X1 port map( A1 => n4675, A2 => n554, B1 => n4707, B2 => n557,
                           ZN => n1839);
   U1895 : NAND4_X1 port map( A1 => n1840, A2 => n1841, A3 => n1842, A4 => 
                           n1843, ZN => n1830);
   U1896 : AOI221_X1 port map( B1 => n560, B2 => n4995, C1 => n563, C2 => n5027
                           , A => n1844, ZN => n1843);
   U1897 : OAI22_X1 port map( A1 => n1845, A2 => n566, B1 => n1846, B2 => n569,
                           ZN => n1844);
   U1898 : AOI221_X1 port map( B1 => n572, B2 => n5283, C1 => n575, C2 => n5251
                           , A => n1847, ZN => n1842);
   U1899 : OAI22_X1 port map( A1 => n1848, A2 => n578, B1 => n1849, B2 => n581,
                           ZN => n1847);
   U1900 : AOI221_X1 port map( B1 => n584, B2 => n4547, C1 => n587, C2 => n4579
                           , A => n1850, ZN => n1841);
   U1901 : OAI22_X1 port map( A1 => n1851, A2 => n590, B1 => n1852, B2 => n593,
                           ZN => n1850);
   U1902 : AOI221_X1 port map( B1 => n596, B2 => n4611, C1 => n599, C2 => n4643
                           , A => n1853, ZN => n1840);
   U1903 : OAI22_X1 port map( A1 => n1854, A2 => n602, B1 => n1855, B2 => n605,
                           ZN => n1853);
   U1904 : MUX2_X1 port map( A => n1856, B => n338, S => n503, Z => n3076);
   U1905 : INV_X1 port map( A => n1857, ZN => n785);
   U1906 : OAI221_X1 port map( B1 => n1857, B2 => n506, C1 => n273, C2 => n1858
                           , A => n1859, ZN => n3075);
   U1907 : OAI21_X1 port map( B1 => n1860, B2 => n1861, A => n509, ZN => n1859)
                           ;
   U1908 : NAND4_X1 port map( A1 => n1862, A2 => n1863, A3 => n1864, A4 => 
                           n1865, ZN => n1861);
   U1909 : AOI221_X1 port map( B1 => n512, B2 => n1047, C1 => n515, C2 => n1013
                           , A => n1866, ZN => n1865);
   U1910 : OAI22_X1 port map( A1 => n5058, A2 => n518, B1 => n5090, B2 => n521,
                           ZN => n1866);
   U1911 : AOI221_X1 port map( B1 => n524, B2 => n875, C1 => n527, C2 => n909, 
                           A => n1867, ZN => n1864);
   U1912 : OAI22_X1 port map( A1 => n5346, A2 => n530, B1 => n5314, B2 => n533,
                           ZN => n1867);
   U1913 : AOI221_X1 port map( B1 => n536, B2 => n1856, C1 => n539, C2 => n1296
                           , A => n1868, ZN => n1863);
   U1914 : OAI22_X1 port map( A1 => n4482, A2 => n542, B1 => n4514, B2 => n545,
                           ZN => n1868);
   U1915 : AOI221_X1 port map( B1 => n548, B2 => n1117, C1 => n551, C2 => n1083
                           , A => n1869, ZN => n1862);
   U1916 : OAI22_X1 port map( A1 => n4674, A2 => n554, B1 => n4706, B2 => n557,
                           ZN => n1869);
   U1917 : NAND4_X1 port map( A1 => n1870, A2 => n1871, A3 => n1872, A4 => 
                           n1873, ZN => n1860);
   U1918 : AOI221_X1 port map( B1 => n560, B2 => n4994, C1 => n563, C2 => n5026
                           , A => n1874, ZN => n1873);
   U1919 : OAI22_X1 port map( A1 => n1875, A2 => n566, B1 => n1876, B2 => n569,
                           ZN => n1874);
   U1920 : AOI221_X1 port map( B1 => n572, B2 => n5282, C1 => n575, C2 => n5250
                           , A => n1877, ZN => n1872);
   U1921 : OAI22_X1 port map( A1 => n1878, A2 => n578, B1 => n1879, B2 => n581,
                           ZN => n1877);
   U1922 : AOI221_X1 port map( B1 => n584, B2 => n4546, C1 => n587, C2 => n4578
                           , A => n1880, ZN => n1871);
   U1923 : OAI22_X1 port map( A1 => n1881, A2 => n590, B1 => n1882, B2 => n593,
                           ZN => n1880);
   U1924 : AOI221_X1 port map( B1 => n596, B2 => n4610, C1 => n599, C2 => n4642
                           , A => n1883, ZN => n1870);
   U1925 : OAI22_X1 port map( A1 => n1884, A2 => n602, B1 => n1885, B2 => n605,
                           ZN => n1883);
   U1926 : MUX2_X1 port map( A => n1886, B => n341, S => n503, Z => n3074);
   U1927 : INV_X1 port map( A => n1887, ZN => n787);
   U1928 : OAI221_X1 port map( B1 => n1887, B2 => n506, C1 => n271, C2 => n1888
                           , A => n1889, ZN => n3073);
   U1929 : OAI21_X1 port map( B1 => n1890, B2 => n1891, A => n509, ZN => n1889)
                           ;
   U1930 : NAND4_X1 port map( A1 => n1892, A2 => n1893, A3 => n1894, A4 => 
                           n1895, ZN => n1891);
   U1931 : AOI221_X1 port map( B1 => n512, B2 => n1048, C1 => n515, C2 => n1014
                           , A => n1896, ZN => n1895);
   U1932 : OAI22_X1 port map( A1 => n5057, A2 => n518, B1 => n5089, B2 => n521,
                           ZN => n1896);
   U1933 : AOI221_X1 port map( B1 => n524, B2 => n876, C1 => n527, C2 => n910, 
                           A => n1897, ZN => n1894);
   U1934 : OAI22_X1 port map( A1 => n5345, A2 => n530, B1 => n5313, B2 => n533,
                           ZN => n1897);
   U1935 : AOI221_X1 port map( B1 => n536, B2 => n1886, C1 => n539, C2 => n1297
                           , A => n1898, ZN => n1893);
   U1936 : OAI22_X1 port map( A1 => n4481, A2 => n542, B1 => n4513, B2 => n545,
                           ZN => n1898);
   U1937 : AOI221_X1 port map( B1 => n548, B2 => n1118, C1 => n551, C2 => n1084
                           , A => n1899, ZN => n1892);
   U1938 : OAI22_X1 port map( A1 => n4673, A2 => n554, B1 => n4705, B2 => n557,
                           ZN => n1899);
   U1939 : NAND4_X1 port map( A1 => n1900, A2 => n1901, A3 => n1902, A4 => 
                           n1903, ZN => n1890);
   U1940 : AOI221_X1 port map( B1 => n560, B2 => n4993, C1 => n563, C2 => n5025
                           , A => n1904, ZN => n1903);
   U1941 : OAI22_X1 port map( A1 => n1905, A2 => n566, B1 => n1906, B2 => n569,
                           ZN => n1904);
   U1942 : AOI221_X1 port map( B1 => n572, B2 => n5281, C1 => n575, C2 => n5249
                           , A => n1907, ZN => n1902);
   U1943 : OAI22_X1 port map( A1 => n1908, A2 => n578, B1 => n1909, B2 => n581,
                           ZN => n1907);
   U1944 : AOI221_X1 port map( B1 => n584, B2 => n4545, C1 => n587, C2 => n4577
                           , A => n1910, ZN => n1901);
   U1945 : OAI22_X1 port map( A1 => n1911, A2 => n590, B1 => n1912, B2 => n593,
                           ZN => n1910);
   U1946 : AOI221_X1 port map( B1 => n596, B2 => n4609, C1 => n599, C2 => n4641
                           , A => n1913, ZN => n1900);
   U1947 : OAI22_X1 port map( A1 => n1914, A2 => n602, B1 => n1915, B2 => n605,
                           ZN => n1913);
   U1948 : MUX2_X1 port map( A => n1916, B => n344, S => n503, Z => n3072);
   U1949 : INV_X1 port map( A => n1917, ZN => n789);
   U1950 : OAI221_X1 port map( B1 => n1917, B2 => n506, C1 => n271, C2 => n1918
                           , A => n1919, ZN => n3071);
   U1951 : OAI21_X1 port map( B1 => n1920, B2 => n1921, A => n509, ZN => n1919)
                           ;
   U1952 : NAND4_X1 port map( A1 => n1922, A2 => n1923, A3 => n1924, A4 => 
                           n1925, ZN => n1921);
   U1953 : AOI221_X1 port map( B1 => n512, B2 => n1049, C1 => n515, C2 => n1015
                           , A => n1926, ZN => n1925);
   U1954 : OAI22_X1 port map( A1 => n5056, A2 => n518, B1 => n5088, B2 => n521,
                           ZN => n1926);
   U1955 : AOI221_X1 port map( B1 => n524, B2 => n877, C1 => n527, C2 => n911, 
                           A => n1927, ZN => n1924);
   U1956 : OAI22_X1 port map( A1 => n5344, A2 => n530, B1 => n5312, B2 => n533,
                           ZN => n1927);
   U1957 : AOI221_X1 port map( B1 => n536, B2 => n1916, C1 => n539, C2 => n1298
                           , A => n1928, ZN => n1923);
   U1958 : OAI22_X1 port map( A1 => n4480, A2 => n542, B1 => n4512, B2 => n545,
                           ZN => n1928);
   U1959 : AOI221_X1 port map( B1 => n548, B2 => n1119, C1 => n551, C2 => n1085
                           , A => n1929, ZN => n1922);
   U1960 : OAI22_X1 port map( A1 => n4672, A2 => n554, B1 => n4704, B2 => n557,
                           ZN => n1929);
   U1961 : NAND4_X1 port map( A1 => n1930, A2 => n1931, A3 => n1932, A4 => 
                           n1933, ZN => n1920);
   U1962 : AOI221_X1 port map( B1 => n560, B2 => n4992, C1 => n563, C2 => n5024
                           , A => n1934, ZN => n1933);
   U1963 : OAI22_X1 port map( A1 => n1935, A2 => n566, B1 => n1936, B2 => n569,
                           ZN => n1934);
   U1964 : AOI221_X1 port map( B1 => n572, B2 => n5280, C1 => n575, C2 => n5248
                           , A => n1937, ZN => n1932);
   U1965 : OAI22_X1 port map( A1 => n1938, A2 => n578, B1 => n1939, B2 => n581,
                           ZN => n1937);
   U1966 : AOI221_X1 port map( B1 => n584, B2 => n4544, C1 => n587, C2 => n4576
                           , A => n1940, ZN => n1931);
   U1967 : OAI22_X1 port map( A1 => n1941, A2 => n590, B1 => n1942, B2 => n593,
                           ZN => n1940);
   U1968 : AOI221_X1 port map( B1 => n596, B2 => n4608, C1 => n599, C2 => n4640
                           , A => n1943, ZN => n1930);
   U1969 : OAI22_X1 port map( A1 => n1944, A2 => n602, B1 => n1945, B2 => n605,
                           ZN => n1943);
   U1970 : MUX2_X1 port map( A => n1946, B => n347, S => n502, Z => n3070);
   U1971 : INV_X1 port map( A => n1947, ZN => n791);
   U1972 : OAI221_X1 port map( B1 => n1947, B2 => n506, C1 => n274, C2 => n1948
                           , A => n1949, ZN => n3069);
   U1973 : OAI21_X1 port map( B1 => n1950, B2 => n1951, A => n508, ZN => n1949)
                           ;
   U1974 : NAND4_X1 port map( A1 => n1952, A2 => n1953, A3 => n1954, A4 => 
                           n1955, ZN => n1951);
   U1975 : AOI221_X1 port map( B1 => n511, B2 => n1050, C1 => n514, C2 => n1016
                           , A => n1956, ZN => n1955);
   U1976 : OAI22_X1 port map( A1 => n5055, A2 => n517, B1 => n5087, B2 => n520,
                           ZN => n1956);
   U1977 : AOI221_X1 port map( B1 => n523, B2 => n878, C1 => n526, C2 => n912, 
                           A => n1957, ZN => n1954);
   U1978 : OAI22_X1 port map( A1 => n5343, A2 => n529, B1 => n5311, B2 => n532,
                           ZN => n1957);
   U1979 : AOI221_X1 port map( B1 => n535, B2 => n1946, C1 => n538, C2 => n1299
                           , A => n1958, ZN => n1953);
   U1980 : OAI22_X1 port map( A1 => n4479, A2 => n541, B1 => n4511, B2 => n544,
                           ZN => n1958);
   U1981 : AOI221_X1 port map( B1 => n547, B2 => n1120, C1 => n550, C2 => n1086
                           , A => n1959, ZN => n1952);
   U1982 : OAI22_X1 port map( A1 => n4671, A2 => n553, B1 => n4703, B2 => n556,
                           ZN => n1959);
   U1983 : NAND4_X1 port map( A1 => n1960, A2 => n1961, A3 => n1962, A4 => 
                           n1963, ZN => n1950);
   U1984 : AOI221_X1 port map( B1 => n559, B2 => n4991, C1 => n562, C2 => n5023
                           , A => n1964, ZN => n1963);
   U1985 : OAI22_X1 port map( A1 => n1965, A2 => n565, B1 => n1966, B2 => n568,
                           ZN => n1964);
   U1986 : AOI221_X1 port map( B1 => n571, B2 => n5279, C1 => n574, C2 => n5247
                           , A => n1967, ZN => n1962);
   U1987 : OAI22_X1 port map( A1 => n1968, A2 => n577, B1 => n1969, B2 => n580,
                           ZN => n1967);
   U1988 : AOI221_X1 port map( B1 => n583, B2 => n4543, C1 => n586, C2 => n4575
                           , A => n1970, ZN => n1961);
   U1989 : OAI22_X1 port map( A1 => n1971, A2 => n589, B1 => n1972, B2 => n592,
                           ZN => n1970);
   U1990 : AOI221_X1 port map( B1 => n595, B2 => n4607, C1 => n598, C2 => n4639
                           , A => n1973, ZN => n1960);
   U1991 : OAI22_X1 port map( A1 => n1974, A2 => n601, B1 => n1975, B2 => n604,
                           ZN => n1973);
   U1992 : MUX2_X1 port map( A => n1976, B => n350, S => n502, Z => n3068);
   U1993 : INV_X1 port map( A => n1977, ZN => n793);
   U1994 : OAI221_X1 port map( B1 => n1977, B2 => n506, C1 => n271, C2 => n1978
                           , A => n1979, ZN => n3067);
   U1995 : OAI21_X1 port map( B1 => n1980, B2 => n1981, A => n508, ZN => n1979)
                           ;
   U1996 : NAND4_X1 port map( A1 => n1982, A2 => n1983, A3 => n1984, A4 => 
                           n1985, ZN => n1981);
   U1997 : AOI221_X1 port map( B1 => n511, B2 => n1051, C1 => n514, C2 => n1017
                           , A => n1986, ZN => n1985);
   U1998 : OAI22_X1 port map( A1 => n5054, A2 => n517, B1 => n5086, B2 => n520,
                           ZN => n1986);
   U1999 : AOI221_X1 port map( B1 => n523, B2 => n879, C1 => n526, C2 => n913, 
                           A => n1987, ZN => n1984);
   U2000 : OAI22_X1 port map( A1 => n5342, A2 => n529, B1 => n5310, B2 => n532,
                           ZN => n1987);
   U2001 : AOI221_X1 port map( B1 => n535, B2 => n1976, C1 => n538, C2 => n1300
                           , A => n1988, ZN => n1983);
   U2002 : OAI22_X1 port map( A1 => n4478, A2 => n541, B1 => n4510, B2 => n544,
                           ZN => n1988);
   U2003 : AOI221_X1 port map( B1 => n547, B2 => n1121, C1 => n550, C2 => n1087
                           , A => n1989, ZN => n1982);
   U2004 : OAI22_X1 port map( A1 => n4670, A2 => n553, B1 => n4702, B2 => n556,
                           ZN => n1989);
   U2005 : NAND4_X1 port map( A1 => n1990, A2 => n1991, A3 => n1992, A4 => 
                           n1993, ZN => n1980);
   U2006 : AOI221_X1 port map( B1 => n559, B2 => n4990, C1 => n562, C2 => n5022
                           , A => n1994, ZN => n1993);
   U2007 : OAI22_X1 port map( A1 => n1995, A2 => n565, B1 => n1996, B2 => n568,
                           ZN => n1994);
   U2008 : AOI221_X1 port map( B1 => n571, B2 => n5278, C1 => n574, C2 => n5246
                           , A => n1997, ZN => n1992);
   U2009 : OAI22_X1 port map( A1 => n1998, A2 => n577, B1 => n1999, B2 => n580,
                           ZN => n1997);
   U2010 : AOI221_X1 port map( B1 => n583, B2 => n4542, C1 => n586, C2 => n4574
                           , A => n2000, ZN => n1991);
   U2011 : OAI22_X1 port map( A1 => n2001, A2 => n589, B1 => n2002, B2 => n592,
                           ZN => n2000);
   U2012 : AOI221_X1 port map( B1 => n595, B2 => n4606, C1 => n598, C2 => n4638
                           , A => n2003, ZN => n1990);
   U2013 : OAI22_X1 port map( A1 => n2004, A2 => n601, B1 => n2005, B2 => n604,
                           ZN => n2003);
   U2014 : MUX2_X1 port map( A => n2006, B => n353, S => n502, Z => n3066);
   U2015 : INV_X1 port map( A => n2007, ZN => n795);
   U2016 : OAI221_X1 port map( B1 => n2007, B2 => n506, C1 => n271, C2 => n2008
                           , A => n2009, ZN => n3065);
   U2017 : OAI21_X1 port map( B1 => n2010, B2 => n2011, A => n508, ZN => n2009)
                           ;
   U2018 : NAND4_X1 port map( A1 => n2012, A2 => n2013, A3 => n2014, A4 => 
                           n2015, ZN => n2011);
   U2019 : AOI221_X1 port map( B1 => n511, B2 => n1052, C1 => n514, C2 => n1018
                           , A => n2016, ZN => n2015);
   U2020 : OAI22_X1 port map( A1 => n5053, A2 => n517, B1 => n5085, B2 => n520,
                           ZN => n2016);
   U2021 : AOI221_X1 port map( B1 => n523, B2 => n880, C1 => n526, C2 => n914, 
                           A => n2017, ZN => n2014);
   U2022 : OAI22_X1 port map( A1 => n5341, A2 => n529, B1 => n5309, B2 => n532,
                           ZN => n2017);
   U2023 : AOI221_X1 port map( B1 => n535, B2 => n2006, C1 => n538, C2 => n1301
                           , A => n2018, ZN => n2013);
   U2024 : OAI22_X1 port map( A1 => n4477, A2 => n541, B1 => n4509, B2 => n544,
                           ZN => n2018);
   U2025 : AOI221_X1 port map( B1 => n547, B2 => n1122, C1 => n550, C2 => n1088
                           , A => n2019, ZN => n2012);
   U2026 : OAI22_X1 port map( A1 => n4669, A2 => n553, B1 => n4701, B2 => n556,
                           ZN => n2019);
   U2027 : NAND4_X1 port map( A1 => n2020, A2 => n2021, A3 => n2022, A4 => 
                           n2023, ZN => n2010);
   U2028 : AOI221_X1 port map( B1 => n559, B2 => n4989, C1 => n562, C2 => n5021
                           , A => n2024, ZN => n2023);
   U2029 : OAI22_X1 port map( A1 => n2025, A2 => n565, B1 => n2026, B2 => n568,
                           ZN => n2024);
   U2030 : AOI221_X1 port map( B1 => n571, B2 => n5277, C1 => n574, C2 => n5245
                           , A => n2027, ZN => n2022);
   U2031 : OAI22_X1 port map( A1 => n2028, A2 => n577, B1 => n2029, B2 => n580,
                           ZN => n2027);
   U2032 : AOI221_X1 port map( B1 => n583, B2 => n4541, C1 => n586, C2 => n4573
                           , A => n2030, ZN => n2021);
   U2033 : OAI22_X1 port map( A1 => n2031, A2 => n589, B1 => n2032, B2 => n592,
                           ZN => n2030);
   U2034 : AOI221_X1 port map( B1 => n595, B2 => n4605, C1 => n598, C2 => n4637
                           , A => n2033, ZN => n2020);
   U2035 : OAI22_X1 port map( A1 => n2034, A2 => n601, B1 => n2035, B2 => n604,
                           ZN => n2033);
   U2036 : MUX2_X1 port map( A => n2036, B => n356, S => n502, Z => n3064);
   U2037 : INV_X1 port map( A => n2037, ZN => n797);
   U2038 : OAI221_X1 port map( B1 => n2037, B2 => n506, C1 => n271, C2 => n2038
                           , A => n2039, ZN => n3063);
   U2039 : OAI21_X1 port map( B1 => n2040, B2 => n2041, A => n508, ZN => n2039)
                           ;
   U2040 : NAND4_X1 port map( A1 => n2042, A2 => n2043, A3 => n2044, A4 => 
                           n2045, ZN => n2041);
   U2041 : AOI221_X1 port map( B1 => n511, B2 => n1053, C1 => n514, C2 => n1019
                           , A => n2046, ZN => n2045);
   U2042 : OAI22_X1 port map( A1 => n5052, A2 => n517, B1 => n5084, B2 => n520,
                           ZN => n2046);
   U2043 : AOI221_X1 port map( B1 => n523, B2 => n881, C1 => n526, C2 => n915, 
                           A => n2047, ZN => n2044);
   U2044 : OAI22_X1 port map( A1 => n5340, A2 => n529, B1 => n5308, B2 => n532,
                           ZN => n2047);
   U2045 : AOI221_X1 port map( B1 => n535, B2 => n2036, C1 => n538, C2 => n1302
                           , A => n2048, ZN => n2043);
   U2046 : OAI22_X1 port map( A1 => n4476, A2 => n541, B1 => n4508, B2 => n544,
                           ZN => n2048);
   U2047 : AOI221_X1 port map( B1 => n547, B2 => n1123, C1 => n550, C2 => n1089
                           , A => n2049, ZN => n2042);
   U2048 : OAI22_X1 port map( A1 => n4668, A2 => n553, B1 => n4700, B2 => n556,
                           ZN => n2049);
   U2049 : NAND4_X1 port map( A1 => n2050, A2 => n2051, A3 => n2052, A4 => 
                           n2053, ZN => n2040);
   U2050 : AOI221_X1 port map( B1 => n559, B2 => n4988, C1 => n562, C2 => n5020
                           , A => n2054, ZN => n2053);
   U2051 : OAI22_X1 port map( A1 => n2055, A2 => n565, B1 => n2056, B2 => n568,
                           ZN => n2054);
   U2052 : AOI221_X1 port map( B1 => n571, B2 => n5276, C1 => n574, C2 => n5244
                           , A => n2057, ZN => n2052);
   U2053 : OAI22_X1 port map( A1 => n2058, A2 => n577, B1 => n2059, B2 => n580,
                           ZN => n2057);
   U2054 : AOI221_X1 port map( B1 => n583, B2 => n4540, C1 => n586, C2 => n4572
                           , A => n2060, ZN => n2051);
   U2055 : OAI22_X1 port map( A1 => n2061, A2 => n589, B1 => n2062, B2 => n592,
                           ZN => n2060);
   U2056 : AOI221_X1 port map( B1 => n595, B2 => n4604, C1 => n598, C2 => n4636
                           , A => n2063, ZN => n2050);
   U2057 : OAI22_X1 port map( A1 => n2064, A2 => n601, B1 => n2065, B2 => n604,
                           ZN => n2063);
   U2058 : MUX2_X1 port map( A => n2066, B => n359, S => n502, Z => n3062);
   U2059 : INV_X1 port map( A => n2067, ZN => n799);
   U2060 : OAI221_X1 port map( B1 => n2067, B2 => n507, C1 => n275, C2 => n2068
                           , A => n2069, ZN => n3061);
   U2061 : OAI21_X1 port map( B1 => n2070, B2 => n2071, A => n508, ZN => n2069)
                           ;
   U2062 : NAND4_X1 port map( A1 => n2072, A2 => n2073, A3 => n2074, A4 => 
                           n2075, ZN => n2071);
   U2063 : AOI221_X1 port map( B1 => n511, B2 => n1054, C1 => n514, C2 => n1020
                           , A => n2076, ZN => n2075);
   U2064 : OAI22_X1 port map( A1 => n5051, A2 => n517, B1 => n5083, B2 => n520,
                           ZN => n2076);
   U2065 : AOI221_X1 port map( B1 => n523, B2 => n882, C1 => n526, C2 => n916, 
                           A => n2077, ZN => n2074);
   U2066 : OAI22_X1 port map( A1 => n5339, A2 => n529, B1 => n5307, B2 => n532,
                           ZN => n2077);
   U2067 : AOI221_X1 port map( B1 => n535, B2 => n2066, C1 => n538, C2 => n1303
                           , A => n2078, ZN => n2073);
   U2068 : OAI22_X1 port map( A1 => n4475, A2 => n541, B1 => n4507, B2 => n544,
                           ZN => n2078);
   U2069 : AOI221_X1 port map( B1 => n547, B2 => n1124, C1 => n550, C2 => n1090
                           , A => n2079, ZN => n2072);
   U2070 : OAI22_X1 port map( A1 => n4667, A2 => n553, B1 => n4699, B2 => n556,
                           ZN => n2079);
   U2071 : NAND4_X1 port map( A1 => n2080, A2 => n2081, A3 => n2082, A4 => 
                           n2083, ZN => n2070);
   U2072 : AOI221_X1 port map( B1 => n559, B2 => n4987, C1 => n562, C2 => n5019
                           , A => n2084, ZN => n2083);
   U2073 : OAI22_X1 port map( A1 => n2085, A2 => n565, B1 => n2086, B2 => n568,
                           ZN => n2084);
   U2074 : AOI221_X1 port map( B1 => n571, B2 => n5275, C1 => n574, C2 => n5243
                           , A => n2087, ZN => n2082);
   U2075 : OAI22_X1 port map( A1 => n2088, A2 => n577, B1 => n2089, B2 => n580,
                           ZN => n2087);
   U2076 : AOI221_X1 port map( B1 => n583, B2 => n4539, C1 => n586, C2 => n4571
                           , A => n2090, ZN => n2081);
   U2077 : OAI22_X1 port map( A1 => n2091, A2 => n589, B1 => n2092, B2 => n592,
                           ZN => n2090);
   U2078 : AOI221_X1 port map( B1 => n595, B2 => n4603, C1 => n598, C2 => n4635
                           , A => n2093, ZN => n2080);
   U2079 : OAI22_X1 port map( A1 => n2094, A2 => n601, B1 => n2095, B2 => n604,
                           ZN => n2093);
   U2080 : MUX2_X1 port map( A => n2096, B => n362, S => n502, Z => n3060);
   U2081 : INV_X1 port map( A => n2097, ZN => n801);
   U2082 : OAI221_X1 port map( B1 => n2097, B2 => n507, C1 => n271, C2 => n2098
                           , A => n2099, ZN => n3059);
   U2083 : OAI21_X1 port map( B1 => n2100, B2 => n2101, A => n508, ZN => n2099)
                           ;
   U2084 : NAND4_X1 port map( A1 => n2102, A2 => n2103, A3 => n2104, A4 => 
                           n2105, ZN => n2101);
   U2085 : AOI221_X1 port map( B1 => n511, B2 => n1055, C1 => n514, C2 => n1021
                           , A => n2106, ZN => n2105);
   U2086 : OAI22_X1 port map( A1 => n5050, A2 => n517, B1 => n5082, B2 => n520,
                           ZN => n2106);
   U2087 : AOI221_X1 port map( B1 => n523, B2 => n883, C1 => n526, C2 => n917, 
                           A => n2107, ZN => n2104);
   U2088 : OAI22_X1 port map( A1 => n5338, A2 => n529, B1 => n5306, B2 => n532,
                           ZN => n2107);
   U2089 : AOI221_X1 port map( B1 => n535, B2 => n2096, C1 => n538, C2 => n1304
                           , A => n2108, ZN => n2103);
   U2090 : OAI22_X1 port map( A1 => n4474, A2 => n541, B1 => n4506, B2 => n544,
                           ZN => n2108);
   U2091 : AOI221_X1 port map( B1 => n547, B2 => n1125, C1 => n550, C2 => n1091
                           , A => n2109, ZN => n2102);
   U2092 : OAI22_X1 port map( A1 => n4666, A2 => n553, B1 => n4698, B2 => n556,
                           ZN => n2109);
   U2093 : NAND4_X1 port map( A1 => n2110, A2 => n2111, A3 => n2112, A4 => 
                           n2113, ZN => n2100);
   U2094 : AOI221_X1 port map( B1 => n559, B2 => n4986, C1 => n562, C2 => n5018
                           , A => n2114, ZN => n2113);
   U2095 : OAI22_X1 port map( A1 => n2115, A2 => n565, B1 => n2116, B2 => n568,
                           ZN => n2114);
   U2096 : AOI221_X1 port map( B1 => n571, B2 => n5274, C1 => n574, C2 => n5242
                           , A => n2117, ZN => n2112);
   U2097 : OAI22_X1 port map( A1 => n2118, A2 => n577, B1 => n2119, B2 => n580,
                           ZN => n2117);
   U2098 : AOI221_X1 port map( B1 => n583, B2 => n4538, C1 => n586, C2 => n4570
                           , A => n2120, ZN => n2111);
   U2099 : OAI22_X1 port map( A1 => n2121, A2 => n589, B1 => n2122, B2 => n592,
                           ZN => n2120);
   U2100 : AOI221_X1 port map( B1 => n595, B2 => n4602, C1 => n598, C2 => n4634
                           , A => n2123, ZN => n2110);
   U2101 : OAI22_X1 port map( A1 => n2124, A2 => n601, B1 => n2125, B2 => n604,
                           ZN => n2123);
   U2102 : MUX2_X1 port map( A => n2126, B => n365, S => n502, Z => n3058);
   U2103 : INV_X1 port map( A => n2127, ZN => n803);
   U2104 : OAI221_X1 port map( B1 => n2127, B2 => n507, C1 => n272, C2 => n2128
                           , A => n2129, ZN => n3057);
   U2105 : OAI21_X1 port map( B1 => n2130, B2 => n2131, A => n508, ZN => n2129)
                           ;
   U2106 : NAND4_X1 port map( A1 => n2132, A2 => n2133, A3 => n2134, A4 => 
                           n2135, ZN => n2131);
   U2107 : AOI221_X1 port map( B1 => n511, B2 => n1056, C1 => n514, C2 => n1022
                           , A => n2136, ZN => n2135);
   U2108 : OAI22_X1 port map( A1 => n5049, A2 => n517, B1 => n5081, B2 => n520,
                           ZN => n2136);
   U2109 : AOI221_X1 port map( B1 => n523, B2 => n884, C1 => n526, C2 => n918, 
                           A => n2137, ZN => n2134);
   U2110 : OAI22_X1 port map( A1 => n5337, A2 => n529, B1 => n5305, B2 => n532,
                           ZN => n2137);
   U2111 : AOI221_X1 port map( B1 => n535, B2 => n2126, C1 => n538, C2 => n1305
                           , A => n2138, ZN => n2133);
   U2112 : OAI22_X1 port map( A1 => n4473, A2 => n541, B1 => n4505, B2 => n544,
                           ZN => n2138);
   U2113 : AOI221_X1 port map( B1 => n547, B2 => n1126, C1 => n550, C2 => n1092
                           , A => n2139, ZN => n2132);
   U2114 : OAI22_X1 port map( A1 => n4665, A2 => n553, B1 => n4697, B2 => n556,
                           ZN => n2139);
   U2115 : NAND4_X1 port map( A1 => n2140, A2 => n2141, A3 => n2142, A4 => 
                           n2143, ZN => n2130);
   U2116 : AOI221_X1 port map( B1 => n559, B2 => n4985, C1 => n562, C2 => n5017
                           , A => n2144, ZN => n2143);
   U2117 : OAI22_X1 port map( A1 => n2145, A2 => n565, B1 => n2146, B2 => n568,
                           ZN => n2144);
   U2118 : AOI221_X1 port map( B1 => n571, B2 => n5273, C1 => n574, C2 => n5241
                           , A => n2147, ZN => n2142);
   U2119 : OAI22_X1 port map( A1 => n2148, A2 => n577, B1 => n2149, B2 => n580,
                           ZN => n2147);
   U2120 : AOI221_X1 port map( B1 => n583, B2 => n4537, C1 => n586, C2 => n4569
                           , A => n2150, ZN => n2141);
   U2121 : OAI22_X1 port map( A1 => n2151, A2 => n589, B1 => n2152, B2 => n592,
                           ZN => n2150);
   U2122 : AOI221_X1 port map( B1 => n595, B2 => n4601, C1 => n598, C2 => n4633
                           , A => n2153, ZN => n2140);
   U2123 : OAI22_X1 port map( A1 => n2154, A2 => n601, B1 => n2155, B2 => n604,
                           ZN => n2153);
   U2124 : MUX2_X1 port map( A => n2156, B => n368, S => n502, Z => n3056);
   U2125 : INV_X1 port map( A => n2157, ZN => n805);
   U2126 : OAI221_X1 port map( B1 => n2157, B2 => n507, C1 => n271, C2 => n2158
                           , A => n2159, ZN => n3055);
   U2127 : OAI21_X1 port map( B1 => n2160, B2 => n2161, A => n508, ZN => n2159)
                           ;
   U2128 : NAND4_X1 port map( A1 => n2162, A2 => n2163, A3 => n2164, A4 => 
                           n2165, ZN => n2161);
   U2129 : AOI221_X1 port map( B1 => n511, B2 => n1057, C1 => n514, C2 => n1023
                           , A => n2166, ZN => n2165);
   U2130 : OAI22_X1 port map( A1 => n5048, A2 => n517, B1 => n5080, B2 => n520,
                           ZN => n2166);
   U2131 : AOI221_X1 port map( B1 => n523, B2 => n885, C1 => n526, C2 => n919, 
                           A => n2167, ZN => n2164);
   U2132 : OAI22_X1 port map( A1 => n5336, A2 => n529, B1 => n5304, B2 => n532,
                           ZN => n2167);
   U2133 : AOI221_X1 port map( B1 => n535, B2 => n2156, C1 => n538, C2 => n1306
                           , A => n2168, ZN => n2163);
   U2134 : OAI22_X1 port map( A1 => n4472, A2 => n541, B1 => n4504, B2 => n544,
                           ZN => n2168);
   U2135 : AOI221_X1 port map( B1 => n547, B2 => n1127, C1 => n550, C2 => n1093
                           , A => n2169, ZN => n2162);
   U2136 : OAI22_X1 port map( A1 => n4664, A2 => n553, B1 => n4696, B2 => n556,
                           ZN => n2169);
   U2137 : NAND4_X1 port map( A1 => n2170, A2 => n2171, A3 => n2172, A4 => 
                           n2173, ZN => n2160);
   U2138 : AOI221_X1 port map( B1 => n559, B2 => n4984, C1 => n562, C2 => n5016
                           , A => n2174, ZN => n2173);
   U2139 : OAI22_X1 port map( A1 => n2175, A2 => n565, B1 => n2176, B2 => n568,
                           ZN => n2174);
   U2140 : AOI221_X1 port map( B1 => n571, B2 => n5272, C1 => n574, C2 => n5240
                           , A => n2177, ZN => n2172);
   U2141 : OAI22_X1 port map( A1 => n2178, A2 => n577, B1 => n2179, B2 => n580,
                           ZN => n2177);
   U2142 : AOI221_X1 port map( B1 => n583, B2 => n4536, C1 => n586, C2 => n4568
                           , A => n2180, ZN => n2171);
   U2143 : OAI22_X1 port map( A1 => n2181, A2 => n589, B1 => n2182, B2 => n592,
                           ZN => n2180);
   U2144 : AOI221_X1 port map( B1 => n595, B2 => n4600, C1 => n598, C2 => n4632
                           , A => n2183, ZN => n2170);
   U2145 : OAI22_X1 port map( A1 => n2184, A2 => n601, B1 => n2185, B2 => n604,
                           ZN => n2183);
   U2146 : MUX2_X1 port map( A => n2186, B => n371, S => n502, Z => n3054);
   U2147 : INV_X1 port map( A => n2187, ZN => n807);
   U2148 : OAI221_X1 port map( B1 => n2187, B2 => n507, C1 => n274, C2 => n2188
                           , A => n2189, ZN => n3053);
   U2149 : OAI21_X1 port map( B1 => n2190, B2 => n2191, A => n508, ZN => n2189)
                           ;
   U2150 : NAND4_X1 port map( A1 => n2192, A2 => n2193, A3 => n2194, A4 => 
                           n2195, ZN => n2191);
   U2151 : AOI221_X1 port map( B1 => n511, B2 => n1058, C1 => n514, C2 => n1024
                           , A => n2196, ZN => n2195);
   U2152 : OAI22_X1 port map( A1 => n5047, A2 => n517, B1 => n5079, B2 => n520,
                           ZN => n2196);
   U2153 : AOI221_X1 port map( B1 => n523, B2 => n886, C1 => n526, C2 => n920, 
                           A => n2197, ZN => n2194);
   U2154 : OAI22_X1 port map( A1 => n5335, A2 => n529, B1 => n5303, B2 => n532,
                           ZN => n2197);
   U2155 : AOI221_X1 port map( B1 => n535, B2 => n2186, C1 => n538, C2 => n1307
                           , A => n2198, ZN => n2193);
   U2156 : OAI22_X1 port map( A1 => n4471, A2 => n541, B1 => n4503, B2 => n544,
                           ZN => n2198);
   U2157 : AOI221_X1 port map( B1 => n547, B2 => n1128, C1 => n550, C2 => n1094
                           , A => n2199, ZN => n2192);
   U2158 : OAI22_X1 port map( A1 => n4663, A2 => n553, B1 => n4695, B2 => n556,
                           ZN => n2199);
   U2159 : NAND4_X1 port map( A1 => n2200, A2 => n2201, A3 => n2202, A4 => 
                           n2203, ZN => n2190);
   U2160 : AOI221_X1 port map( B1 => n559, B2 => n4983, C1 => n562, C2 => n5015
                           , A => n2204, ZN => n2203);
   U2161 : OAI22_X1 port map( A1 => n2205, A2 => n565, B1 => n2206, B2 => n568,
                           ZN => n2204);
   U2162 : AOI221_X1 port map( B1 => n571, B2 => n5271, C1 => n574, C2 => n5239
                           , A => n2207, ZN => n2202);
   U2163 : OAI22_X1 port map( A1 => n2208, A2 => n577, B1 => n2209, B2 => n580,
                           ZN => n2207);
   U2164 : AOI221_X1 port map( B1 => n583, B2 => n4535, C1 => n586, C2 => n4567
                           , A => n2210, ZN => n2201);
   U2165 : OAI22_X1 port map( A1 => n2211, A2 => n589, B1 => n2212, B2 => n592,
                           ZN => n2210);
   U2166 : AOI221_X1 port map( B1 => n595, B2 => n4599, C1 => n598, C2 => n4631
                           , A => n2213, ZN => n2200);
   U2167 : OAI22_X1 port map( A1 => n2214, A2 => n601, B1 => n2215, B2 => n604,
                           ZN => n2213);
   U2168 : MUX2_X1 port map( A => n2216, B => n374, S => n502, Z => n3052);
   U2169 : INV_X1 port map( A => n2217, ZN => n809);
   U2170 : OAI221_X1 port map( B1 => n2217, B2 => n507, C1 => n270, C2 => n2218
                           , A => n2219, ZN => n3051);
   U2171 : OAI21_X1 port map( B1 => n2220, B2 => n2221, A => n508, ZN => n2219)
                           ;
   U2172 : NAND4_X1 port map( A1 => n2222, A2 => n2223, A3 => n2224, A4 => 
                           n2225, ZN => n2221);
   U2173 : AOI221_X1 port map( B1 => n511, B2 => n1059, C1 => n514, C2 => n1025
                           , A => n2226, ZN => n2225);
   U2174 : OAI22_X1 port map( A1 => n5046, A2 => n517, B1 => n5078, B2 => n520,
                           ZN => n2226);
   U2175 : AOI221_X1 port map( B1 => n523, B2 => n887, C1 => n526, C2 => n921, 
                           A => n2227, ZN => n2224);
   U2176 : OAI22_X1 port map( A1 => n5334, A2 => n529, B1 => n5302, B2 => n532,
                           ZN => n2227);
   U2177 : AOI221_X1 port map( B1 => n535, B2 => n2216, C1 => n538, C2 => n1308
                           , A => n2228, ZN => n2223);
   U2178 : OAI22_X1 port map( A1 => n4470, A2 => n541, B1 => n4502, B2 => n544,
                           ZN => n2228);
   U2179 : AOI221_X1 port map( B1 => n547, B2 => n1129, C1 => n550, C2 => n1095
                           , A => n2229, ZN => n2222);
   U2180 : OAI22_X1 port map( A1 => n4662, A2 => n553, B1 => n4694, B2 => n556,
                           ZN => n2229);
   U2181 : NAND4_X1 port map( A1 => n2230, A2 => n2231, A3 => n2232, A4 => 
                           n2233, ZN => n2220);
   U2182 : AOI221_X1 port map( B1 => n559, B2 => n4982, C1 => n562, C2 => n5014
                           , A => n2234, ZN => n2233);
   U2183 : OAI22_X1 port map( A1 => n2235, A2 => n565, B1 => n2236, B2 => n568,
                           ZN => n2234);
   U2184 : AOI221_X1 port map( B1 => n571, B2 => n5270, C1 => n574, C2 => n5238
                           , A => n2237, ZN => n2232);
   U2185 : OAI22_X1 port map( A1 => n2238, A2 => n577, B1 => n2239, B2 => n580,
                           ZN => n2237);
   U2186 : AOI221_X1 port map( B1 => n583, B2 => n4534, C1 => n586, C2 => n4566
                           , A => n2240, ZN => n2231);
   U2187 : OAI22_X1 port map( A1 => n2241, A2 => n589, B1 => n2242, B2 => n592,
                           ZN => n2240);
   U2188 : AOI221_X1 port map( B1 => n595, B2 => n4598, C1 => n598, C2 => n4630
                           , A => n2243, ZN => n2230);
   U2189 : OAI22_X1 port map( A1 => n2244, A2 => n601, B1 => n2245, B2 => n604,
                           ZN => n2243);
   U2190 : MUX2_X1 port map( A => n2246, B => n377, S => n502, Z => n3050);
   U2191 : INV_X1 port map( A => n2247, ZN => n811);
   U2192 : OAI221_X1 port map( B1 => n2247, B2 => n507, C1 => n270, C2 => n2248
                           , A => n2249, ZN => n3049);
   U2193 : OAI21_X1 port map( B1 => n2250, B2 => n2251, A => n508, ZN => n2249)
                           ;
   U2194 : NAND4_X1 port map( A1 => n2252, A2 => n2253, A3 => n2254, A4 => 
                           n2255, ZN => n2251);
   U2195 : AOI221_X1 port map( B1 => n511, B2 => n1060, C1 => n514, C2 => n1026
                           , A => n2256, ZN => n2255);
   U2196 : OAI22_X1 port map( A1 => n5045, A2 => n517, B1 => n5077, B2 => n520,
                           ZN => n2256);
   U2197 : AOI221_X1 port map( B1 => n523, B2 => n888, C1 => n526, C2 => n922, 
                           A => n2257, ZN => n2254);
   U2198 : OAI22_X1 port map( A1 => n5333, A2 => n529, B1 => n5301, B2 => n532,
                           ZN => n2257);
   U2199 : AOI221_X1 port map( B1 => n535, B2 => n2246, C1 => n538, C2 => n1309
                           , A => n2258, ZN => n2253);
   U2200 : OAI22_X1 port map( A1 => n4469, A2 => n541, B1 => n4501, B2 => n544,
                           ZN => n2258);
   U2201 : AOI221_X1 port map( B1 => n547, B2 => n1130, C1 => n550, C2 => n1096
                           , A => n2259, ZN => n2252);
   U2202 : OAI22_X1 port map( A1 => n4661, A2 => n553, B1 => n4693, B2 => n556,
                           ZN => n2259);
   U2203 : NAND4_X1 port map( A1 => n2260, A2 => n2261, A3 => n2262, A4 => 
                           n2263, ZN => n2250);
   U2204 : AOI221_X1 port map( B1 => n559, B2 => n4981, C1 => n562, C2 => n5013
                           , A => n2264, ZN => n2263);
   U2205 : OAI22_X1 port map( A1 => n2265, A2 => n565, B1 => n2266, B2 => n568,
                           ZN => n2264);
   U2206 : AOI221_X1 port map( B1 => n571, B2 => n5269, C1 => n574, C2 => n5237
                           , A => n2267, ZN => n2262);
   U2207 : OAI22_X1 port map( A1 => n2268, A2 => n577, B1 => n2269, B2 => n580,
                           ZN => n2267);
   U2208 : AOI221_X1 port map( B1 => n583, B2 => n4533, C1 => n586, C2 => n4565
                           , A => n2270, ZN => n2261);
   U2209 : OAI22_X1 port map( A1 => n2271, A2 => n589, B1 => n2272, B2 => n592,
                           ZN => n2270);
   U2210 : AOI221_X1 port map( B1 => n595, B2 => n4597, C1 => n598, C2 => n4629
                           , A => n2273, ZN => n2260);
   U2211 : OAI22_X1 port map( A1 => n2274, A2 => n601, B1 => n2275, B2 => n604,
                           ZN => n2273);
   U2212 : MUX2_X1 port map( A => n2276, B => n380, S => n502, Z => n3048);
   U2213 : OAI21_X1 port map( B1 => n853, B2 => n1274, A => n260, ZN => n1312);
   U2214 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => ADD_WR(2), A3 => n1134, ZN
                           => n1274);
   U2215 : AND3_X1 port map( A1 => WR, A2 => ENABLE, A3 => ADD_WR(4), ZN => 
                           n1134);
   U2216 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), ZN => n853);
   U2217 : INV_X1 port map( A => n2277, ZN => n813);
   U2218 : OAI221_X1 port map( B1 => n2277, B2 => n507, C1 => n273, C2 => n2278
                           , A => n2279, ZN => n3047);
   U2219 : OAI21_X1 port map( B1 => n2280, B2 => n2281, A => n508, ZN => n2279)
                           ;
   U2220 : AND2_X1 port map( A1 => n507, A2 => n276, ZN => n1319);
   U2221 : NAND4_X1 port map( A1 => n2282, A2 => n2283, A3 => n2284, A4 => 
                           n2285, ZN => n2281);
   U2222 : AOI221_X1 port map( B1 => n511, B2 => n1061, C1 => n514, C2 => n1027
                           , A => n2286, ZN => n2285);
   U2223 : OAI22_X1 port map( A1 => n5044, A2 => n517, B1 => n5076, B2 => n520,
                           ZN => n2286);
   U2224 : NAND2_X1 port map( A1 => n2287, A2 => n2288, ZN => n1328);
   U2225 : NAND2_X1 port map( A1 => n2287, A2 => n2289, ZN => n1327);
   U2226 : AND2_X1 port map( A1 => n2290, A2 => n2288, ZN => n1325);
   U2227 : AND2_X1 port map( A1 => n2290, A2 => n2289, ZN => n1324);
   U2228 : AOI221_X1 port map( B1 => n523, B2 => n889, C1 => n526, C2 => n923, 
                           A => n2291, ZN => n2284);
   U2229 : OAI22_X1 port map( A1 => n5332, A2 => n529, B1 => n5300, B2 => n532,
                           ZN => n2291);
   U2230 : NAND2_X1 port map( A1 => n2287, A2 => n2292, ZN => n1333);
   U2231 : NAND2_X1 port map( A1 => n2287, A2 => n2293, ZN => n1332);
   U2232 : AND2_X1 port map( A1 => n2290, A2 => n2292, ZN => n1330);
   U2233 : AND2_X1 port map( A1 => n2290, A2 => n2293, ZN => n1329);
   U2234 : AOI221_X1 port map( B1 => n535, B2 => n2276, C1 => n538, C2 => n1310
                           , A => n2294, ZN => n2283);
   U2235 : OAI22_X1 port map( A1 => n4468, A2 => n541, B1 => n4500, B2 => n544,
                           ZN => n2294);
   U2236 : NAND2_X1 port map( A1 => n2295, A2 => n2296, ZN => n1338);
   U2237 : NAND2_X1 port map( A1 => n2297, A2 => n2296, ZN => n1337);
   U2238 : AND2_X1 port map( A1 => n2295, A2 => n2298, ZN => n1335);
   U2239 : AND2_X1 port map( A1 => n2297, A2 => n2298, ZN => n1334);
   U2240 : AOI221_X1 port map( B1 => n547, B2 => n1131, C1 => n550, C2 => n1097
                           , A => n2299, ZN => n2282);
   U2241 : OAI22_X1 port map( A1 => n4660, A2 => n553, B1 => n4692, B2 => n556,
                           ZN => n2299);
   U2242 : NAND2_X1 port map( A1 => n2300, A2 => n2290, ZN => n1343);
   U2243 : NAND2_X1 port map( A1 => n2301, A2 => n2290, ZN => n1342);
   U2244 : AND2_X1 port map( A1 => n2300, A2 => n2287, ZN => n1340);
   U2245 : AND2_X1 port map( A1 => n2301, A2 => n2287, ZN => n1339);
   U2246 : NAND4_X1 port map( A1 => n2302, A2 => n2303, A3 => n2304, A4 => 
                           n2305, ZN => n2280);
   U2247 : AOI221_X1 port map( B1 => n559, B2 => n4980, C1 => n562, C2 => n5012
                           , A => n2306, ZN => n2305);
   U2248 : OAI22_X1 port map( A1 => n2307, A2 => n565, B1 => n2308, B2 => n568,
                           ZN => n2306);
   U2249 : NAND2_X1 port map( A1 => n2298, A2 => n2288, ZN => n1354);
   U2250 : NAND2_X1 port map( A1 => n2298, A2 => n2289, ZN => n1352);
   U2251 : AND2_X1 port map( A1 => n2288, A2 => n2296, ZN => n1349);
   U2252 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(4), A3 => n2309, 
                           ZN => n2288);
   U2253 : AND2_X1 port map( A1 => n2296, A2 => n2289, ZN => n1348);
   U2254 : NOR3_X1 port map( A1 => n2310, A2 => ADD_RD2(4), A3 => n2309, ZN => 
                           n2289);
   U2255 : AOI221_X1 port map( B1 => n571, B2 => n5268, C1 => n574, C2 => n5236
                           , A => n2311, ZN => n2304);
   U2256 : OAI22_X1 port map( A1 => n2312, A2 => n577, B1 => n2313, B2 => n580,
                           ZN => n2311);
   U2257 : NAND2_X1 port map( A1 => n2292, A2 => n2298, ZN => n1361);
   U2258 : NAND2_X1 port map( A1 => n2293, A2 => n2298, ZN => n1359);
   U2259 : AND2_X1 port map( A1 => n2292, A2 => n2296, ZN => n1356);
   U2260 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => n2310, 
                           ZN => n2292);
   U2261 : AND2_X1 port map( A1 => n2293, A2 => n2296, ZN => n1355);
   U2262 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => 
                           ADD_RD2(0), ZN => n2293);
   U2263 : AOI221_X1 port map( B1 => n583, B2 => n4532, C1 => n586, C2 => n4564
                           , A => n2314, ZN => n2303);
   U2264 : OAI22_X1 port map( A1 => n2315, A2 => n589, B1 => n2316, B2 => n592,
                           ZN => n2314);
   U2265 : NAND2_X1 port map( A1 => n2290, A2 => n2295, ZN => n1368);
   U2266 : NAND2_X1 port map( A1 => n2290, A2 => n2297, ZN => n1366);
   U2267 : NOR2_X1 port map( A1 => n2317, A2 => ADD_RD2(1), ZN => n2290);
   U2268 : AND2_X1 port map( A1 => n2295, A2 => n2287, ZN => n1363);
   U2269 : NOR3_X1 port map( A1 => n2318, A2 => ADD_RD2(0), A3 => n2309, ZN => 
                           n2295);
   U2270 : AND2_X1 port map( A1 => n2287, A2 => n2297, ZN => n1362);
   U2271 : NOR3_X1 port map( A1 => n2318, A2 => n2310, A3 => n2309, ZN => n2297
                           );
   U2272 : NOR2_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), ZN => n2287);
   U2273 : AOI221_X1 port map( B1 => n595, B2 => n4596, C1 => n598, C2 => n4628
                           , A => n2319, ZN => n2302);
   U2274 : OAI22_X1 port map( A1 => n2320, A2 => n601, B1 => n2321, B2 => n604,
                           ZN => n2319);
   U2275 : NAND2_X1 port map( A1 => n2300, A2 => n2296, ZN => n1375);
   U2276 : NAND2_X1 port map( A1 => n2301, A2 => n2296, ZN => n1373);
   U2277 : NOR2_X1 port map( A1 => n2322, A2 => ADD_RD2(2), ZN => n2296);
   U2278 : AND2_X1 port map( A1 => n2300, A2 => n2298, ZN => n1370);
   U2279 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(3), A3 => n2318, 
                           ZN => n2300);
   U2280 : AND2_X1 port map( A1 => n2301, A2 => n2298, ZN => n1369);
   U2281 : NOR2_X1 port map( A1 => n2317, A2 => n2322, ZN => n2298);
   U2282 : INV_X1 port map( A => ADD_RD2(1), ZN => n2322);
   U2283 : NOR3_X1 port map( A1 => n2310, A2 => ADD_RD2(3), A3 => n2318, ZN => 
                           n2301);
   U2284 : INV_X1 port map( A => ADD_RD2(0), ZN => n2310);
   U2285 : NAND4_X1 port map( A1 => n2323, A2 => n2324, A3 => n2325, A4 => 
                           n2326, ZN => n1314);
   U2286 : NOR4_X1 port map( A1 => n748, A2 => n1064, A3 => n2327, A4 => n2328,
                           ZN => n2326);
   U2287 : XOR2_X1 port map( A => ADD_WR(1), B => ADD_RD2(1), Z => n2328);
   U2288 : XOR2_X1 port map( A => ADD_WR(0), B => ADD_RD2(0), Z => n2327);
   U2289 : INV_X1 port map( A => RD2, ZN => n748);
   U2290 : XOR2_X1 port map( A => n2309, B => ADD_WR(3), Z => n2325);
   U2291 : INV_X1 port map( A => ADD_RD2(3), ZN => n2309);
   U2292 : XOR2_X1 port map( A => ADD_WR(4), B => n2318, Z => n2324);
   U2293 : INV_X1 port map( A => ADD_RD2(4), ZN => n2318);
   U2294 : XOR2_X1 port map( A => n2317, B => ADD_WR(2), Z => n2323);
   U2295 : INV_X1 port map( A => ADD_RD2(2), ZN => n2317);
   U2296 : OAI221_X1 port map( B1 => n1313, B2 => n607, C1 => n275, C2 => n2330
                           , A => n2331, ZN => n3046);
   U2297 : OAI21_X1 port map( B1 => n2332, B2 => n2333, A => n612, ZN => n2331)
                           ;
   U2298 : NAND4_X1 port map( A1 => n2335, A2 => n2336, A3 => n2337, A4 => 
                           n2338, ZN => n2333);
   U2299 : AOI221_X1 port map( B1 => n615, B2 => n1029, C1 => n618, C2 => n995,
                           A => n2341, ZN => n2338);
   U2300 : OAI22_X1 port map( A1 => n5075, A2 => n621, B1 => n5107, B2 => n624,
                           ZN => n2341);
   U2301 : AOI221_X1 port map( B1 => n627, B2 => n857, C1 => n630, C2 => n891, 
                           A => n2346, ZN => n2337);
   U2302 : OAI22_X1 port map( A1 => n5363, A2 => n633, B1 => n5331, B2 => n636,
                           ZN => n2346);
   U2303 : AOI221_X1 port map( B1 => n639, B2 => n1311, C1 => n642, C2 => n1278
                           , A => n2351, ZN => n2336);
   U2304 : OAI22_X1 port map( A1 => n4499, A2 => n645, B1 => n4531, B2 => n648,
                           ZN => n2351);
   U2305 : AOI221_X1 port map( B1 => n651, B2 => n1099, C1 => n654, C2 => n1065
                           , A => n2356, ZN => n2335);
   U2306 : OAI22_X1 port map( A1 => n4691, A2 => n657, B1 => n4723, B2 => n660,
                           ZN => n2356);
   U2307 : NAND4_X1 port map( A1 => n2359, A2 => n2360, A3 => n2361, A4 => 
                           n2362, ZN => n2332);
   U2308 : AOI221_X1 port map( B1 => n663, B2 => n5011, C1 => n666, C2 => n5043
                           , A => n2365, ZN => n2362);
   U2309 : OAI22_X1 port map( A1 => n1351, A2 => n669, B1 => n1353, B2 => n672,
                           ZN => n2365);
   U2310 : AOI221_X1 port map( B1 => n675, B2 => n5299, C1 => n678, C2 => n5267
                           , A => n2370, ZN => n2361);
   U2311 : OAI22_X1 port map( A1 => n1358, A2 => n681, B1 => n1360, B2 => n684,
                           ZN => n2370);
   U2312 : AOI221_X1 port map( B1 => n687, B2 => n4563, C1 => n690, C2 => n4595
                           , A => n2375, ZN => n2360);
   U2313 : OAI22_X1 port map( A1 => n1365, A2 => n693, B1 => n1367, B2 => n696,
                           ZN => n2375);
   U2314 : AOI221_X1 port map( B1 => n699, B2 => n4627, C1 => n702, C2 => n4659
                           , A => n2380, ZN => n2359);
   U2315 : OAI22_X1 port map( A1 => n1372, A2 => n705, B1 => n1374, B2 => n708,
                           ZN => n2380);
   U2316 : NAND2_X1 port map( A1 => DATAIN(31), A2 => n265, ZN => n1313);
   U2317 : OAI21_X1 port map( B1 => n269, B2 => n2383, A => n712, ZN => n3045);
   U2318 : OAI221_X1 port map( B1 => n1377, B2 => n607, C1 => n272, C2 => n2385
                           , A => n2386, ZN => n3044);
   U2319 : OAI21_X1 port map( B1 => n2387, B2 => n2388, A => n612, ZN => n2386)
                           ;
   U2320 : NAND4_X1 port map( A1 => n2389, A2 => n2390, A3 => n2391, A4 => 
                           n2392, ZN => n2388);
   U2321 : AOI221_X1 port map( B1 => n615, B2 => n1031, C1 => n618, C2 => n997,
                           A => n2393, ZN => n2392);
   U2322 : OAI22_X1 port map( A1 => n5074, A2 => n621, B1 => n5106, B2 => n624,
                           ZN => n2393);
   U2323 : AOI221_X1 port map( B1 => n627, B2 => n859, C1 => n630, C2 => n893, 
                           A => n2394, ZN => n2391);
   U2324 : OAI22_X1 port map( A1 => n5362, A2 => n633, B1 => n5330, B2 => n636,
                           ZN => n2394);
   U2325 : AOI221_X1 port map( B1 => n639, B2 => n1376, C1 => n642, C2 => n1280
                           , A => n2395, ZN => n2390);
   U2326 : OAI22_X1 port map( A1 => n4498, A2 => n645, B1 => n4530, B2 => n648,
                           ZN => n2395);
   U2327 : AOI221_X1 port map( B1 => n651, B2 => n1101, C1 => n654, C2 => n1067
                           , A => n2396, ZN => n2389);
   U2328 : OAI22_X1 port map( A1 => n4690, A2 => n657, B1 => n4722, B2 => n660,
                           ZN => n2396);
   U2329 : NAND4_X1 port map( A1 => n2397, A2 => n2398, A3 => n2399, A4 => 
                           n2400, ZN => n2387);
   U2330 : AOI221_X1 port map( B1 => n663, B2 => n5010, C1 => n666, C2 => n5042
                           , A => n2401, ZN => n2400);
   U2331 : OAI22_X1 port map( A1 => n1395, A2 => n669, B1 => n1396, B2 => n672,
                           ZN => n2401);
   U2332 : AOI221_X1 port map( B1 => n675, B2 => n5298, C1 => n678, C2 => n5266
                           , A => n2402, ZN => n2399);
   U2333 : OAI22_X1 port map( A1 => n1398, A2 => n681, B1 => n1399, B2 => n684,
                           ZN => n2402);
   U2334 : AOI221_X1 port map( B1 => n687, B2 => n4562, C1 => n690, C2 => n4594
                           , A => n2403, ZN => n2398);
   U2335 : OAI22_X1 port map( A1 => n1401, A2 => n693, B1 => n1402, B2 => n696,
                           ZN => n2403);
   U2336 : AOI221_X1 port map( B1 => n699, B2 => n4626, C1 => n702, C2 => n4658
                           , A => n2404, ZN => n2397);
   U2337 : OAI22_X1 port map( A1 => n1404, A2 => n705, B1 => n1405, B2 => n708,
                           ZN => n2404);
   U2338 : NAND2_X1 port map( A1 => DATAIN(30), A2 => n264, ZN => n1377);
   U2339 : OAI21_X1 port map( B1 => n268, B2 => n2405, A => n712, ZN => n3043);
   U2340 : OAI221_X1 port map( B1 => n1407, B2 => n607, C1 => n272, C2 => n2406
                           , A => n2407, ZN => n3042);
   U2341 : OAI21_X1 port map( B1 => n2408, B2 => n2409, A => n612, ZN => n2407)
                           ;
   U2342 : NAND4_X1 port map( A1 => n2410, A2 => n2411, A3 => n2412, A4 => 
                           n2413, ZN => n2409);
   U2343 : AOI221_X1 port map( B1 => n615, B2 => n1032, C1 => n618, C2 => n998,
                           A => n2414, ZN => n2413);
   U2344 : OAI22_X1 port map( A1 => n5073, A2 => n621, B1 => n5105, B2 => n624,
                           ZN => n2414);
   U2345 : AOI221_X1 port map( B1 => n627, B2 => n860, C1 => n630, C2 => n894, 
                           A => n2415, ZN => n2412);
   U2346 : OAI22_X1 port map( A1 => n5361, A2 => n633, B1 => n5329, B2 => n636,
                           ZN => n2415);
   U2347 : AOI221_X1 port map( B1 => n639, B2 => n1406, C1 => n642, C2 => n1281
                           , A => n2416, ZN => n2411);
   U2348 : OAI22_X1 port map( A1 => n4497, A2 => n645, B1 => n4529, B2 => n648,
                           ZN => n2416);
   U2349 : AOI221_X1 port map( B1 => n651, B2 => n1102, C1 => n654, C2 => n1068
                           , A => n2417, ZN => n2410);
   U2350 : OAI22_X1 port map( A1 => n4689, A2 => n657, B1 => n4721, B2 => n660,
                           ZN => n2417);
   U2351 : NAND4_X1 port map( A1 => n2418, A2 => n2419, A3 => n2420, A4 => 
                           n2421, ZN => n2408);
   U2352 : AOI221_X1 port map( B1 => n663, B2 => n5009, C1 => n666, C2 => n5041
                           , A => n2422, ZN => n2421);
   U2353 : OAI22_X1 port map( A1 => n1425, A2 => n669, B1 => n1426, B2 => n672,
                           ZN => n2422);
   U2354 : AOI221_X1 port map( B1 => n675, B2 => n5297, C1 => n678, C2 => n5265
                           , A => n2423, ZN => n2420);
   U2355 : OAI22_X1 port map( A1 => n1428, A2 => n681, B1 => n1429, B2 => n684,
                           ZN => n2423);
   U2356 : AOI221_X1 port map( B1 => n687, B2 => n4561, C1 => n690, C2 => n4593
                           , A => n2424, ZN => n2419);
   U2357 : OAI22_X1 port map( A1 => n1431, A2 => n693, B1 => n1432, B2 => n696,
                           ZN => n2424);
   U2358 : AOI221_X1 port map( B1 => n699, B2 => n4625, C1 => n702, C2 => n4657
                           , A => n2425, ZN => n2418);
   U2359 : OAI22_X1 port map( A1 => n1434, A2 => n705, B1 => n1435, B2 => n708,
                           ZN => n2425);
   U2360 : NAND2_X1 port map( A1 => DATAIN(29), A2 => n265, ZN => n1407);
   U2361 : OAI21_X1 port map( B1 => n269, B2 => n2426, A => n712, ZN => n3041);
   U2362 : OAI221_X1 port map( B1 => n1437, B2 => n607, C1 => n272, C2 => n2427
                           , A => n2428, ZN => n3040);
   U2363 : OAI21_X1 port map( B1 => n2429, B2 => n2430, A => n612, ZN => n2428)
                           ;
   U2364 : NAND4_X1 port map( A1 => n2431, A2 => n2432, A3 => n2433, A4 => 
                           n2434, ZN => n2430);
   U2365 : AOI221_X1 port map( B1 => n615, B2 => n1033, C1 => n618, C2 => n999,
                           A => n2435, ZN => n2434);
   U2366 : OAI22_X1 port map( A1 => n5072, A2 => n621, B1 => n5104, B2 => n624,
                           ZN => n2435);
   U2367 : AOI221_X1 port map( B1 => n627, B2 => n861, C1 => n630, C2 => n895, 
                           A => n2436, ZN => n2433);
   U2368 : OAI22_X1 port map( A1 => n5360, A2 => n633, B1 => n5328, B2 => n636,
                           ZN => n2436);
   U2369 : AOI221_X1 port map( B1 => n639, B2 => n1436, C1 => n642, C2 => n1282
                           , A => n2437, ZN => n2432);
   U2370 : OAI22_X1 port map( A1 => n4496, A2 => n645, B1 => n4528, B2 => n648,
                           ZN => n2437);
   U2371 : AOI221_X1 port map( B1 => n651, B2 => n1103, C1 => n654, C2 => n1069
                           , A => n2438, ZN => n2431);
   U2372 : OAI22_X1 port map( A1 => n4688, A2 => n657, B1 => n4720, B2 => n660,
                           ZN => n2438);
   U2373 : NAND4_X1 port map( A1 => n2439, A2 => n2440, A3 => n2441, A4 => 
                           n2442, ZN => n2429);
   U2374 : AOI221_X1 port map( B1 => n663, B2 => n5008, C1 => n666, C2 => n5040
                           , A => n2443, ZN => n2442);
   U2375 : OAI22_X1 port map( A1 => n1455, A2 => n669, B1 => n1456, B2 => n672,
                           ZN => n2443);
   U2376 : AOI221_X1 port map( B1 => n675, B2 => n5296, C1 => n678, C2 => n5264
                           , A => n2444, ZN => n2441);
   U2377 : OAI22_X1 port map( A1 => n1458, A2 => n681, B1 => n1459, B2 => n684,
                           ZN => n2444);
   U2378 : AOI221_X1 port map( B1 => n687, B2 => n4560, C1 => n690, C2 => n4592
                           , A => n2445, ZN => n2440);
   U2379 : OAI22_X1 port map( A1 => n1461, A2 => n693, B1 => n1462, B2 => n696,
                           ZN => n2445);
   U2380 : AOI221_X1 port map( B1 => n699, B2 => n4624, C1 => n702, C2 => n4656
                           , A => n2446, ZN => n2439);
   U2381 : OAI22_X1 port map( A1 => n1464, A2 => n705, B1 => n1465, B2 => n708,
                           ZN => n2446);
   U2382 : NAND2_X1 port map( A1 => DATAIN(28), A2 => n265, ZN => n1437);
   U2383 : OAI21_X1 port map( B1 => n268, B2 => n2447, A => n712, ZN => n3039);
   U2384 : OAI221_X1 port map( B1 => n1467, B2 => n607, C1 => n272, C2 => n2448
                           , A => n2449, ZN => n3038);
   U2385 : OAI21_X1 port map( B1 => n2450, B2 => n2451, A => n612, ZN => n2449)
                           ;
   U2386 : NAND4_X1 port map( A1 => n2452, A2 => n2453, A3 => n2454, A4 => 
                           n2455, ZN => n2451);
   U2387 : AOI221_X1 port map( B1 => n615, B2 => n1034, C1 => n618, C2 => n1000
                           , A => n2456, ZN => n2455);
   U2388 : OAI22_X1 port map( A1 => n5071, A2 => n621, B1 => n5103, B2 => n624,
                           ZN => n2456);
   U2389 : AOI221_X1 port map( B1 => n627, B2 => n862, C1 => n630, C2 => n896, 
                           A => n2457, ZN => n2454);
   U2390 : OAI22_X1 port map( A1 => n5359, A2 => n633, B1 => n5327, B2 => n636,
                           ZN => n2457);
   U2391 : AOI221_X1 port map( B1 => n639, B2 => n1466, C1 => n642, C2 => n1283
                           , A => n2458, ZN => n2453);
   U2392 : OAI22_X1 port map( A1 => n4495, A2 => n645, B1 => n4527, B2 => n648,
                           ZN => n2458);
   U2393 : AOI221_X1 port map( B1 => n651, B2 => n1104, C1 => n654, C2 => n1070
                           , A => n2459, ZN => n2452);
   U2394 : OAI22_X1 port map( A1 => n4687, A2 => n657, B1 => n4719, B2 => n660,
                           ZN => n2459);
   U2395 : NAND4_X1 port map( A1 => n2460, A2 => n2461, A3 => n2462, A4 => 
                           n2463, ZN => n2450);
   U2396 : AOI221_X1 port map( B1 => n663, B2 => n5007, C1 => n666, C2 => n5039
                           , A => n2464, ZN => n2463);
   U2397 : OAI22_X1 port map( A1 => n1485, A2 => n669, B1 => n1486, B2 => n672,
                           ZN => n2464);
   U2398 : AOI221_X1 port map( B1 => n675, B2 => n5295, C1 => n678, C2 => n5263
                           , A => n2465, ZN => n2462);
   U2399 : OAI22_X1 port map( A1 => n1488, A2 => n681, B1 => n1489, B2 => n684,
                           ZN => n2465);
   U2400 : AOI221_X1 port map( B1 => n687, B2 => n4559, C1 => n690, C2 => n4591
                           , A => n2466, ZN => n2461);
   U2401 : OAI22_X1 port map( A1 => n1491, A2 => n693, B1 => n1492, B2 => n696,
                           ZN => n2466);
   U2402 : AOI221_X1 port map( B1 => n699, B2 => n4623, C1 => n702, C2 => n4655
                           , A => n2467, ZN => n2460);
   U2403 : OAI22_X1 port map( A1 => n1494, A2 => n705, B1 => n1495, B2 => n708,
                           ZN => n2467);
   U2404 : NAND2_X1 port map( A1 => DATAIN(27), A2 => n265, ZN => n1467);
   U2405 : OAI21_X1 port map( B1 => n268, B2 => n2468, A => n712, ZN => n3037);
   U2406 : OAI221_X1 port map( B1 => n1497, B2 => n607, C1 => n273, C2 => n2469
                           , A => n2470, ZN => n3036);
   U2407 : OAI21_X1 port map( B1 => n2471, B2 => n2472, A => n612, ZN => n2470)
                           ;
   U2408 : NAND4_X1 port map( A1 => n2473, A2 => n2474, A3 => n2475, A4 => 
                           n2476, ZN => n2472);
   U2409 : AOI221_X1 port map( B1 => n615, B2 => n1035, C1 => n618, C2 => n1001
                           , A => n2477, ZN => n2476);
   U2410 : OAI22_X1 port map( A1 => n5070, A2 => n621, B1 => n5102, B2 => n624,
                           ZN => n2477);
   U2411 : AOI221_X1 port map( B1 => n627, B2 => n863, C1 => n630, C2 => n897, 
                           A => n2478, ZN => n2475);
   U2412 : OAI22_X1 port map( A1 => n5358, A2 => n633, B1 => n5326, B2 => n636,
                           ZN => n2478);
   U2413 : AOI221_X1 port map( B1 => n639, B2 => n1496, C1 => n642, C2 => n1284
                           , A => n2479, ZN => n2474);
   U2414 : OAI22_X1 port map( A1 => n4494, A2 => n645, B1 => n4526, B2 => n648,
                           ZN => n2479);
   U2415 : AOI221_X1 port map( B1 => n651, B2 => n1105, C1 => n654, C2 => n1071
                           , A => n2480, ZN => n2473);
   U2416 : OAI22_X1 port map( A1 => n4686, A2 => n657, B1 => n4718, B2 => n660,
                           ZN => n2480);
   U2417 : NAND4_X1 port map( A1 => n2481, A2 => n2482, A3 => n2483, A4 => 
                           n2484, ZN => n2471);
   U2418 : AOI221_X1 port map( B1 => n663, B2 => n5006, C1 => n666, C2 => n5038
                           , A => n2485, ZN => n2484);
   U2419 : OAI22_X1 port map( A1 => n1515, A2 => n669, B1 => n1516, B2 => n672,
                           ZN => n2485);
   U2420 : AOI221_X1 port map( B1 => n675, B2 => n5294, C1 => n678, C2 => n5262
                           , A => n2486, ZN => n2483);
   U2421 : OAI22_X1 port map( A1 => n1518, A2 => n681, B1 => n1519, B2 => n684,
                           ZN => n2486);
   U2422 : AOI221_X1 port map( B1 => n687, B2 => n4558, C1 => n690, C2 => n4590
                           , A => n2487, ZN => n2482);
   U2423 : OAI22_X1 port map( A1 => n1521, A2 => n693, B1 => n1522, B2 => n696,
                           ZN => n2487);
   U2424 : AOI221_X1 port map( B1 => n699, B2 => n4622, C1 => n702, C2 => n4654
                           , A => n2488, ZN => n2481);
   U2425 : OAI22_X1 port map( A1 => n1524, A2 => n705, B1 => n1525, B2 => n708,
                           ZN => n2488);
   U2426 : NAND2_X1 port map( A1 => DATAIN(26), A2 => n264, ZN => n1497);
   U2427 : OAI21_X1 port map( B1 => n268, B2 => n2489, A => n712, ZN => n3035);
   U2428 : OAI221_X1 port map( B1 => n1527, B2 => n607, C1 => n273, C2 => n2490
                           , A => n2491, ZN => n3034);
   U2429 : OAI21_X1 port map( B1 => n2492, B2 => n2493, A => n612, ZN => n2491)
                           ;
   U2430 : NAND4_X1 port map( A1 => n2494, A2 => n2495, A3 => n2496, A4 => 
                           n2497, ZN => n2493);
   U2431 : AOI221_X1 port map( B1 => n615, B2 => n1036, C1 => n618, C2 => n1002
                           , A => n2498, ZN => n2497);
   U2432 : OAI22_X1 port map( A1 => n5069, A2 => n621, B1 => n5101, B2 => n624,
                           ZN => n2498);
   U2433 : AOI221_X1 port map( B1 => n627, B2 => n864, C1 => n630, C2 => n898, 
                           A => n2499, ZN => n2496);
   U2434 : OAI22_X1 port map( A1 => n5357, A2 => n633, B1 => n5325, B2 => n636,
                           ZN => n2499);
   U2435 : AOI221_X1 port map( B1 => n639, B2 => n1526, C1 => n642, C2 => n1285
                           , A => n2500, ZN => n2495);
   U2436 : OAI22_X1 port map( A1 => n4493, A2 => n645, B1 => n4525, B2 => n648,
                           ZN => n2500);
   U2437 : AOI221_X1 port map( B1 => n651, B2 => n1106, C1 => n654, C2 => n1072
                           , A => n2501, ZN => n2494);
   U2438 : OAI22_X1 port map( A1 => n4685, A2 => n657, B1 => n4717, B2 => n660,
                           ZN => n2501);
   U2439 : NAND4_X1 port map( A1 => n2502, A2 => n2503, A3 => n2504, A4 => 
                           n2505, ZN => n2492);
   U2440 : AOI221_X1 port map( B1 => n663, B2 => n5005, C1 => n666, C2 => n5037
                           , A => n2506, ZN => n2505);
   U2441 : OAI22_X1 port map( A1 => n1545, A2 => n669, B1 => n1546, B2 => n672,
                           ZN => n2506);
   U2442 : AOI221_X1 port map( B1 => n675, B2 => n5293, C1 => n678, C2 => n5261
                           , A => n2507, ZN => n2504);
   U2443 : OAI22_X1 port map( A1 => n1548, A2 => n681, B1 => n1549, B2 => n684,
                           ZN => n2507);
   U2444 : AOI221_X1 port map( B1 => n687, B2 => n4557, C1 => n690, C2 => n4589
                           , A => n2508, ZN => n2503);
   U2445 : OAI22_X1 port map( A1 => n1551, A2 => n693, B1 => n1552, B2 => n696,
                           ZN => n2508);
   U2446 : AOI221_X1 port map( B1 => n699, B2 => n4621, C1 => n702, C2 => n4653
                           , A => n2509, ZN => n2502);
   U2447 : OAI22_X1 port map( A1 => n1554, A2 => n705, B1 => n1555, B2 => n708,
                           ZN => n2509);
   U2448 : NAND2_X1 port map( A1 => DATAIN(25), A2 => n265, ZN => n1527);
   U2449 : OAI21_X1 port map( B1 => n269, B2 => n2510, A => n712, ZN => n3033);
   U2450 : OAI221_X1 port map( B1 => n1557, B2 => n607, C1 => n273, C2 => n2511
                           , A => n2512, ZN => n3032);
   U2451 : OAI21_X1 port map( B1 => n2513, B2 => n2514, A => n612, ZN => n2512)
                           ;
   U2452 : NAND4_X1 port map( A1 => n2515, A2 => n2516, A3 => n2517, A4 => 
                           n2518, ZN => n2514);
   U2453 : AOI221_X1 port map( B1 => n615, B2 => n1037, C1 => n618, C2 => n1003
                           , A => n2519, ZN => n2518);
   U2454 : OAI22_X1 port map( A1 => n5068, A2 => n621, B1 => n5100, B2 => n624,
                           ZN => n2519);
   U2455 : AOI221_X1 port map( B1 => n627, B2 => n865, C1 => n630, C2 => n899, 
                           A => n2520, ZN => n2517);
   U2456 : OAI22_X1 port map( A1 => n5356, A2 => n633, B1 => n5324, B2 => n636,
                           ZN => n2520);
   U2457 : AOI221_X1 port map( B1 => n639, B2 => n1556, C1 => n642, C2 => n1286
                           , A => n2521, ZN => n2516);
   U2458 : OAI22_X1 port map( A1 => n4492, A2 => n645, B1 => n4524, B2 => n648,
                           ZN => n2521);
   U2459 : AOI221_X1 port map( B1 => n651, B2 => n1107, C1 => n654, C2 => n1073
                           , A => n2522, ZN => n2515);
   U2460 : OAI22_X1 port map( A1 => n4684, A2 => n657, B1 => n4716, B2 => n660,
                           ZN => n2522);
   U2461 : NAND4_X1 port map( A1 => n2523, A2 => n2524, A3 => n2525, A4 => 
                           n2526, ZN => n2513);
   U2462 : AOI221_X1 port map( B1 => n663, B2 => n5004, C1 => n666, C2 => n5036
                           , A => n2527, ZN => n2526);
   U2463 : OAI22_X1 port map( A1 => n1575, A2 => n669, B1 => n1576, B2 => n672,
                           ZN => n2527);
   U2464 : AOI221_X1 port map( B1 => n675, B2 => n5292, C1 => n678, C2 => n5260
                           , A => n2528, ZN => n2525);
   U2465 : OAI22_X1 port map( A1 => n1578, A2 => n681, B1 => n1579, B2 => n684,
                           ZN => n2528);
   U2466 : AOI221_X1 port map( B1 => n687, B2 => n4556, C1 => n690, C2 => n4588
                           , A => n2529, ZN => n2524);
   U2467 : OAI22_X1 port map( A1 => n1581, A2 => n693, B1 => n1582, B2 => n696,
                           ZN => n2529);
   U2468 : AOI221_X1 port map( B1 => n699, B2 => n4620, C1 => n702, C2 => n4652
                           , A => n2530, ZN => n2523);
   U2469 : OAI22_X1 port map( A1 => n1584, A2 => n705, B1 => n1585, B2 => n708,
                           ZN => n2530);
   U2470 : NAND2_X1 port map( A1 => DATAIN(24), A2 => n265, ZN => n1557);
   U2471 : OAI21_X1 port map( B1 => n268, B2 => n2531, A => n712, ZN => n3031);
   U2472 : OAI221_X1 port map( B1 => n1587, B2 => n607, C1 => n273, C2 => n2532
                           , A => n2533, ZN => n3030);
   U2473 : OAI21_X1 port map( B1 => n2534, B2 => n2535, A => n611, ZN => n2533)
                           ;
   U2474 : NAND4_X1 port map( A1 => n2536, A2 => n2537, A3 => n2538, A4 => 
                           n2539, ZN => n2535);
   U2475 : AOI221_X1 port map( B1 => n614, B2 => n1038, C1 => n617, C2 => n1004
                           , A => n2540, ZN => n2539);
   U2476 : OAI22_X1 port map( A1 => n5067, A2 => n620, B1 => n5099, B2 => n623,
                           ZN => n2540);
   U2477 : AOI221_X1 port map( B1 => n626, B2 => n866, C1 => n629, C2 => n900, 
                           A => n2541, ZN => n2538);
   U2478 : OAI22_X1 port map( A1 => n5355, A2 => n632, B1 => n5323, B2 => n635,
                           ZN => n2541);
   U2479 : AOI221_X1 port map( B1 => n638, B2 => n1586, C1 => n641, C2 => n1287
                           , A => n2542, ZN => n2537);
   U2480 : OAI22_X1 port map( A1 => n4491, A2 => n644, B1 => n4523, B2 => n647,
                           ZN => n2542);
   U2481 : AOI221_X1 port map( B1 => n650, B2 => n1108, C1 => n653, C2 => n1074
                           , A => n2543, ZN => n2536);
   U2482 : OAI22_X1 port map( A1 => n4683, A2 => n656, B1 => n4715, B2 => n659,
                           ZN => n2543);
   U2483 : NAND4_X1 port map( A1 => n2544, A2 => n2545, A3 => n2546, A4 => 
                           n2547, ZN => n2534);
   U2484 : AOI221_X1 port map( B1 => n662, B2 => n5003, C1 => n665, C2 => n5035
                           , A => n2548, ZN => n2547);
   U2485 : OAI22_X1 port map( A1 => n1605, A2 => n668, B1 => n1606, B2 => n671,
                           ZN => n2548);
   U2486 : AOI221_X1 port map( B1 => n674, B2 => n5291, C1 => n677, C2 => n5259
                           , A => n2549, ZN => n2546);
   U2487 : OAI22_X1 port map( A1 => n1608, A2 => n680, B1 => n1609, B2 => n683,
                           ZN => n2549);
   U2488 : AOI221_X1 port map( B1 => n686, B2 => n4555, C1 => n689, C2 => n4587
                           , A => n2550, ZN => n2545);
   U2489 : OAI22_X1 port map( A1 => n1611, A2 => n692, B1 => n1612, B2 => n695,
                           ZN => n2550);
   U2490 : AOI221_X1 port map( B1 => n698, B2 => n4619, C1 => n701, C2 => n4651
                           , A => n2551, ZN => n2544);
   U2491 : OAI22_X1 port map( A1 => n1614, A2 => n704, B1 => n1615, B2 => n707,
                           ZN => n2551);
   U2492 : NAND2_X1 port map( A1 => DATAIN(23), A2 => n264, ZN => n1587);
   U2493 : OAI21_X1 port map( B1 => n269, B2 => n2552, A => n711, ZN => n3029);
   U2494 : OAI221_X1 port map( B1 => n1617, B2 => n607, C1 => n274, C2 => n2553
                           , A => n2554, ZN => n3028);
   U2495 : OAI21_X1 port map( B1 => n2555, B2 => n2556, A => n611, ZN => n2554)
                           ;
   U2496 : NAND4_X1 port map( A1 => n2557, A2 => n2558, A3 => n2559, A4 => 
                           n2560, ZN => n2556);
   U2497 : AOI221_X1 port map( B1 => n614, B2 => n1039, C1 => n617, C2 => n1005
                           , A => n2561, ZN => n2560);
   U2498 : OAI22_X1 port map( A1 => n5066, A2 => n620, B1 => n5098, B2 => n623,
                           ZN => n2561);
   U2499 : AOI221_X1 port map( B1 => n626, B2 => n867, C1 => n629, C2 => n901, 
                           A => n2562, ZN => n2559);
   U2500 : OAI22_X1 port map( A1 => n5354, A2 => n632, B1 => n5322, B2 => n635,
                           ZN => n2562);
   U2501 : AOI221_X1 port map( B1 => n638, B2 => n1616, C1 => n641, C2 => n1288
                           , A => n2563, ZN => n2558);
   U2502 : OAI22_X1 port map( A1 => n4490, A2 => n644, B1 => n4522, B2 => n647,
                           ZN => n2563);
   U2503 : AOI221_X1 port map( B1 => n650, B2 => n1109, C1 => n653, C2 => n1075
                           , A => n2564, ZN => n2557);
   U2504 : OAI22_X1 port map( A1 => n4682, A2 => n656, B1 => n4714, B2 => n659,
                           ZN => n2564);
   U2505 : NAND4_X1 port map( A1 => n2565, A2 => n2566, A3 => n2567, A4 => 
                           n2568, ZN => n2555);
   U2506 : AOI221_X1 port map( B1 => n662, B2 => n5002, C1 => n665, C2 => n5034
                           , A => n2569, ZN => n2568);
   U2507 : OAI22_X1 port map( A1 => n1635, A2 => n668, B1 => n1636, B2 => n671,
                           ZN => n2569);
   U2508 : AOI221_X1 port map( B1 => n674, B2 => n5290, C1 => n677, C2 => n5258
                           , A => n2570, ZN => n2567);
   U2509 : OAI22_X1 port map( A1 => n1638, A2 => n680, B1 => n1639, B2 => n683,
                           ZN => n2570);
   U2510 : AOI221_X1 port map( B1 => n686, B2 => n4554, C1 => n689, C2 => n4586
                           , A => n2571, ZN => n2566);
   U2511 : OAI22_X1 port map( A1 => n1641, A2 => n692, B1 => n1642, B2 => n695,
                           ZN => n2571);
   U2512 : AOI221_X1 port map( B1 => n698, B2 => n4618, C1 => n701, C2 => n4650
                           , A => n2572, ZN => n2565);
   U2513 : OAI22_X1 port map( A1 => n1644, A2 => n704, B1 => n1645, B2 => n707,
                           ZN => n2572);
   U2514 : NAND2_X1 port map( A1 => DATAIN(22), A2 => n264, ZN => n1617);
   U2515 : OAI21_X1 port map( B1 => n268, B2 => n2573, A => n711, ZN => n3027);
   U2516 : OAI221_X1 port map( B1 => n1647, B2 => n607, C1 => n273, C2 => n2574
                           , A => n2575, ZN => n3026);
   U2517 : OAI21_X1 port map( B1 => n2576, B2 => n2577, A => n611, ZN => n2575)
                           ;
   U2518 : NAND4_X1 port map( A1 => n2578, A2 => n2579, A3 => n2580, A4 => 
                           n2581, ZN => n2577);
   U2519 : AOI221_X1 port map( B1 => n614, B2 => n1040, C1 => n617, C2 => n1006
                           , A => n2582, ZN => n2581);
   U2520 : OAI22_X1 port map( A1 => n5065, A2 => n620, B1 => n5097, B2 => n623,
                           ZN => n2582);
   U2521 : AOI221_X1 port map( B1 => n626, B2 => n868, C1 => n629, C2 => n902, 
                           A => n2583, ZN => n2580);
   U2522 : OAI22_X1 port map( A1 => n5353, A2 => n632, B1 => n5321, B2 => n635,
                           ZN => n2583);
   U2523 : AOI221_X1 port map( B1 => n638, B2 => n1646, C1 => n641, C2 => n1289
                           , A => n2584, ZN => n2579);
   U2524 : OAI22_X1 port map( A1 => n4489, A2 => n644, B1 => n4521, B2 => n647,
                           ZN => n2584);
   U2525 : AOI221_X1 port map( B1 => n650, B2 => n1110, C1 => n653, C2 => n1076
                           , A => n2585, ZN => n2578);
   U2526 : OAI22_X1 port map( A1 => n4681, A2 => n656, B1 => n4713, B2 => n659,
                           ZN => n2585);
   U2527 : NAND4_X1 port map( A1 => n2586, A2 => n2587, A3 => n2588, A4 => 
                           n2589, ZN => n2576);
   U2528 : AOI221_X1 port map( B1 => n662, B2 => n5001, C1 => n665, C2 => n5033
                           , A => n2590, ZN => n2589);
   U2529 : OAI22_X1 port map( A1 => n1665, A2 => n668, B1 => n1666, B2 => n671,
                           ZN => n2590);
   U2530 : AOI221_X1 port map( B1 => n674, B2 => n5289, C1 => n677, C2 => n5257
                           , A => n2591, ZN => n2588);
   U2531 : OAI22_X1 port map( A1 => n1668, A2 => n680, B1 => n1669, B2 => n683,
                           ZN => n2591);
   U2532 : AOI221_X1 port map( B1 => n686, B2 => n4553, C1 => n689, C2 => n4585
                           , A => n2592, ZN => n2587);
   U2533 : OAI22_X1 port map( A1 => n1671, A2 => n692, B1 => n1672, B2 => n695,
                           ZN => n2592);
   U2534 : AOI221_X1 port map( B1 => n698, B2 => n4617, C1 => n701, C2 => n4649
                           , A => n2593, ZN => n2586);
   U2535 : OAI22_X1 port map( A1 => n1674, A2 => n704, B1 => n1675, B2 => n707,
                           ZN => n2593);
   U2536 : NAND2_X1 port map( A1 => DATAIN(21), A2 => n264, ZN => n1647);
   U2537 : OAI21_X1 port map( B1 => n269, B2 => n2594, A => n711, ZN => n3025);
   U2538 : OAI221_X1 port map( B1 => n1677, B2 => n607, C1 => n273, C2 => n2595
                           , A => n2596, ZN => n3024);
   U2539 : OAI21_X1 port map( B1 => n2597, B2 => n2598, A => n611, ZN => n2596)
                           ;
   U2540 : NAND4_X1 port map( A1 => n2599, A2 => n2600, A3 => n2601, A4 => 
                           n2602, ZN => n2598);
   U2541 : AOI221_X1 port map( B1 => n614, B2 => n1041, C1 => n617, C2 => n1007
                           , A => n2603, ZN => n2602);
   U2542 : OAI22_X1 port map( A1 => n5064, A2 => n620, B1 => n5096, B2 => n623,
                           ZN => n2603);
   U2543 : AOI221_X1 port map( B1 => n626, B2 => n869, C1 => n629, C2 => n903, 
                           A => n2604, ZN => n2601);
   U2544 : OAI22_X1 port map( A1 => n5352, A2 => n632, B1 => n5320, B2 => n635,
                           ZN => n2604);
   U2545 : AOI221_X1 port map( B1 => n638, B2 => n1676, C1 => n641, C2 => n1290
                           , A => n2605, ZN => n2600);
   U2546 : OAI22_X1 port map( A1 => n4488, A2 => n644, B1 => n4520, B2 => n647,
                           ZN => n2605);
   U2547 : AOI221_X1 port map( B1 => n650, B2 => n1111, C1 => n653, C2 => n1077
                           , A => n2606, ZN => n2599);
   U2548 : OAI22_X1 port map( A1 => n4680, A2 => n656, B1 => n4712, B2 => n659,
                           ZN => n2606);
   U2549 : NAND4_X1 port map( A1 => n2607, A2 => n2608, A3 => n2609, A4 => 
                           n2610, ZN => n2597);
   U2550 : AOI221_X1 port map( B1 => n662, B2 => n5000, C1 => n665, C2 => n5032
                           , A => n2611, ZN => n2610);
   U2551 : OAI22_X1 port map( A1 => n1695, A2 => n668, B1 => n1696, B2 => n671,
                           ZN => n2611);
   U2552 : AOI221_X1 port map( B1 => n674, B2 => n5288, C1 => n677, C2 => n5256
                           , A => n2612, ZN => n2609);
   U2553 : OAI22_X1 port map( A1 => n1698, A2 => n680, B1 => n1699, B2 => n683,
                           ZN => n2612);
   U2554 : AOI221_X1 port map( B1 => n686, B2 => n4552, C1 => n689, C2 => n4584
                           , A => n2613, ZN => n2608);
   U2555 : OAI22_X1 port map( A1 => n1701, A2 => n692, B1 => n1702, B2 => n695,
                           ZN => n2613);
   U2556 : AOI221_X1 port map( B1 => n698, B2 => n4616, C1 => n701, C2 => n4648
                           , A => n2614, ZN => n2607);
   U2557 : OAI22_X1 port map( A1 => n1704, A2 => n704, B1 => n1705, B2 => n707,
                           ZN => n2614);
   U2558 : NAND2_X1 port map( A1 => DATAIN(20), A2 => n264, ZN => n1677);
   U2559 : OAI21_X1 port map( B1 => n268, B2 => n2615, A => n711, ZN => n3023);
   U2560 : OAI221_X1 port map( B1 => n1707, B2 => n608, C1 => n273, C2 => n2616
                           , A => n2617, ZN => n3022);
   U2561 : OAI21_X1 port map( B1 => n2618, B2 => n2619, A => n611, ZN => n2617)
                           ;
   U2562 : NAND4_X1 port map( A1 => n2620, A2 => n2621, A3 => n2622, A4 => 
                           n2623, ZN => n2619);
   U2563 : AOI221_X1 port map( B1 => n614, B2 => n1042, C1 => n617, C2 => n1008
                           , A => n2624, ZN => n2623);
   U2564 : OAI22_X1 port map( A1 => n5063, A2 => n620, B1 => n5095, B2 => n623,
                           ZN => n2624);
   U2565 : AOI221_X1 port map( B1 => n626, B2 => n870, C1 => n629, C2 => n904, 
                           A => n2625, ZN => n2622);
   U2566 : OAI22_X1 port map( A1 => n5351, A2 => n632, B1 => n5319, B2 => n635,
                           ZN => n2625);
   U2567 : AOI221_X1 port map( B1 => n638, B2 => n1706, C1 => n641, C2 => n1291
                           , A => n2626, ZN => n2621);
   U2568 : OAI22_X1 port map( A1 => n4487, A2 => n644, B1 => n4519, B2 => n647,
                           ZN => n2626);
   U2569 : AOI221_X1 port map( B1 => n650, B2 => n1112, C1 => n653, C2 => n1078
                           , A => n2627, ZN => n2620);
   U2570 : OAI22_X1 port map( A1 => n4679, A2 => n656, B1 => n4711, B2 => n659,
                           ZN => n2627);
   U2571 : NAND4_X1 port map( A1 => n2628, A2 => n2629, A3 => n2630, A4 => 
                           n2631, ZN => n2618);
   U2572 : AOI221_X1 port map( B1 => n662, B2 => n4999, C1 => n665, C2 => n5031
                           , A => n2632, ZN => n2631);
   U2573 : OAI22_X1 port map( A1 => n1725, A2 => n668, B1 => n1726, B2 => n671,
                           ZN => n2632);
   U2574 : AOI221_X1 port map( B1 => n674, B2 => n5287, C1 => n677, C2 => n5255
                           , A => n2633, ZN => n2630);
   U2575 : OAI22_X1 port map( A1 => n1728, A2 => n680, B1 => n1729, B2 => n683,
                           ZN => n2633);
   U2576 : AOI221_X1 port map( B1 => n686, B2 => n4551, C1 => n689, C2 => n4583
                           , A => n2634, ZN => n2629);
   U2577 : OAI22_X1 port map( A1 => n1731, A2 => n692, B1 => n1732, B2 => n695,
                           ZN => n2634);
   U2578 : AOI221_X1 port map( B1 => n698, B2 => n4615, C1 => n701, C2 => n4647
                           , A => n2635, ZN => n2628);
   U2579 : OAI22_X1 port map( A1 => n1734, A2 => n704, B1 => n1735, B2 => n707,
                           ZN => n2635);
   U2580 : NAND2_X1 port map( A1 => DATAIN(19), A2 => n264, ZN => n1707);
   U2581 : OAI21_X1 port map( B1 => n270, B2 => n2636, A => n711, ZN => n3021);
   U2582 : OAI221_X1 port map( B1 => n1737, B2 => n608, C1 => n273, C2 => n2637
                           , A => n2638, ZN => n3020);
   U2583 : OAI21_X1 port map( B1 => n2639, B2 => n2640, A => n611, ZN => n2638)
                           ;
   U2584 : NAND4_X1 port map( A1 => n2641, A2 => n2642, A3 => n2643, A4 => 
                           n2644, ZN => n2640);
   U2585 : AOI221_X1 port map( B1 => n614, B2 => n1043, C1 => n617, C2 => n1009
                           , A => n2645, ZN => n2644);
   U2586 : OAI22_X1 port map( A1 => n5062, A2 => n620, B1 => n5094, B2 => n623,
                           ZN => n2645);
   U2587 : AOI221_X1 port map( B1 => n626, B2 => n871, C1 => n629, C2 => n905, 
                           A => n2646, ZN => n2643);
   U2588 : OAI22_X1 port map( A1 => n5350, A2 => n632, B1 => n5318, B2 => n635,
                           ZN => n2646);
   U2589 : AOI221_X1 port map( B1 => n638, B2 => n1736, C1 => n641, C2 => n1292
                           , A => n2647, ZN => n2642);
   U2590 : OAI22_X1 port map( A1 => n4486, A2 => n644, B1 => n4518, B2 => n647,
                           ZN => n2647);
   U2591 : AOI221_X1 port map( B1 => n650, B2 => n1113, C1 => n653, C2 => n1079
                           , A => n2648, ZN => n2641);
   U2592 : OAI22_X1 port map( A1 => n4678, A2 => n656, B1 => n4710, B2 => n659,
                           ZN => n2648);
   U2593 : NAND4_X1 port map( A1 => n2649, A2 => n2650, A3 => n2651, A4 => 
                           n2652, ZN => n2639);
   U2594 : AOI221_X1 port map( B1 => n662, B2 => n4998, C1 => n665, C2 => n5030
                           , A => n2653, ZN => n2652);
   U2595 : OAI22_X1 port map( A1 => n1755, A2 => n668, B1 => n1756, B2 => n671,
                           ZN => n2653);
   U2596 : AOI221_X1 port map( B1 => n674, B2 => n5286, C1 => n677, C2 => n5254
                           , A => n2654, ZN => n2651);
   U2597 : OAI22_X1 port map( A1 => n1758, A2 => n680, B1 => n1759, B2 => n683,
                           ZN => n2654);
   U2598 : AOI221_X1 port map( B1 => n686, B2 => n4550, C1 => n689, C2 => n4582
                           , A => n2655, ZN => n2650);
   U2599 : OAI22_X1 port map( A1 => n1761, A2 => n692, B1 => n1762, B2 => n695,
                           ZN => n2655);
   U2600 : AOI221_X1 port map( B1 => n698, B2 => n4614, C1 => n701, C2 => n4646
                           , A => n2656, ZN => n2649);
   U2601 : OAI22_X1 port map( A1 => n1764, A2 => n704, B1 => n1765, B2 => n707,
                           ZN => n2656);
   U2602 : NAND2_X1 port map( A1 => DATAIN(18), A2 => n263, ZN => n1737);
   U2603 : OAI21_X1 port map( B1 => n268, B2 => n2657, A => n711, ZN => n3019);
   U2604 : OAI221_X1 port map( B1 => n1767, B2 => n608, C1 => n273, C2 => n2658
                           , A => n2659, ZN => n3018);
   U2605 : OAI21_X1 port map( B1 => n2660, B2 => n2661, A => n611, ZN => n2659)
                           ;
   U2606 : NAND4_X1 port map( A1 => n2662, A2 => n2663, A3 => n2664, A4 => 
                           n2665, ZN => n2661);
   U2607 : AOI221_X1 port map( B1 => n614, B2 => n1044, C1 => n617, C2 => n1010
                           , A => n2666, ZN => n2665);
   U2608 : OAI22_X1 port map( A1 => n5061, A2 => n620, B1 => n5093, B2 => n623,
                           ZN => n2666);
   U2609 : AOI221_X1 port map( B1 => n626, B2 => n872, C1 => n629, C2 => n906, 
                           A => n2667, ZN => n2664);
   U2610 : OAI22_X1 port map( A1 => n5349, A2 => n632, B1 => n5317, B2 => n635,
                           ZN => n2667);
   U2611 : AOI221_X1 port map( B1 => n638, B2 => n1766, C1 => n641, C2 => n1293
                           , A => n2668, ZN => n2663);
   U2612 : OAI22_X1 port map( A1 => n4485, A2 => n644, B1 => n4517, B2 => n647,
                           ZN => n2668);
   U2613 : AOI221_X1 port map( B1 => n650, B2 => n1114, C1 => n653, C2 => n1080
                           , A => n2669, ZN => n2662);
   U2614 : OAI22_X1 port map( A1 => n4677, A2 => n656, B1 => n4709, B2 => n659,
                           ZN => n2669);
   U2615 : NAND4_X1 port map( A1 => n2670, A2 => n2671, A3 => n2672, A4 => 
                           n2673, ZN => n2660);
   U2616 : AOI221_X1 port map( B1 => n662, B2 => n4997, C1 => n665, C2 => n5029
                           , A => n2674, ZN => n2673);
   U2617 : OAI22_X1 port map( A1 => n1785, A2 => n668, B1 => n1786, B2 => n671,
                           ZN => n2674);
   U2618 : AOI221_X1 port map( B1 => n674, B2 => n5285, C1 => n677, C2 => n5253
                           , A => n2675, ZN => n2672);
   U2619 : OAI22_X1 port map( A1 => n1788, A2 => n680, B1 => n1789, B2 => n683,
                           ZN => n2675);
   U2620 : AOI221_X1 port map( B1 => n686, B2 => n4549, C1 => n689, C2 => n4581
                           , A => n2676, ZN => n2671);
   U2621 : OAI22_X1 port map( A1 => n1791, A2 => n692, B1 => n1792, B2 => n695,
                           ZN => n2676);
   U2622 : AOI221_X1 port map( B1 => n698, B2 => n4613, C1 => n701, C2 => n4645
                           , A => n2677, ZN => n2670);
   U2623 : OAI22_X1 port map( A1 => n1794, A2 => n704, B1 => n1795, B2 => n707,
                           ZN => n2677);
   U2624 : NAND2_X1 port map( A1 => DATAIN(17), A2 => n264, ZN => n1767);
   U2625 : OAI21_X1 port map( B1 => n270, B2 => n2678, A => n711, ZN => n3017);
   U2626 : OAI221_X1 port map( B1 => n1797, B2 => n608, C1 => n274, C2 => n2679
                           , A => n2680, ZN => n3016);
   U2627 : OAI21_X1 port map( B1 => n2681, B2 => n2682, A => n611, ZN => n2680)
                           ;
   U2628 : NAND4_X1 port map( A1 => n2683, A2 => n2684, A3 => n2685, A4 => 
                           n2686, ZN => n2682);
   U2629 : AOI221_X1 port map( B1 => n614, B2 => n1045, C1 => n617, C2 => n1011
                           , A => n2687, ZN => n2686);
   U2630 : OAI22_X1 port map( A1 => n5060, A2 => n620, B1 => n5092, B2 => n623,
                           ZN => n2687);
   U2631 : AOI221_X1 port map( B1 => n626, B2 => n873, C1 => n629, C2 => n907, 
                           A => n2688, ZN => n2685);
   U2632 : OAI22_X1 port map( A1 => n5348, A2 => n632, B1 => n5316, B2 => n635,
                           ZN => n2688);
   U2633 : AOI221_X1 port map( B1 => n638, B2 => n1796, C1 => n641, C2 => n1294
                           , A => n2689, ZN => n2684);
   U2634 : OAI22_X1 port map( A1 => n4484, A2 => n644, B1 => n4516, B2 => n647,
                           ZN => n2689);
   U2635 : AOI221_X1 port map( B1 => n650, B2 => n1115, C1 => n653, C2 => n1081
                           , A => n2690, ZN => n2683);
   U2636 : OAI22_X1 port map( A1 => n4676, A2 => n656, B1 => n4708, B2 => n659,
                           ZN => n2690);
   U2637 : NAND4_X1 port map( A1 => n2691, A2 => n2692, A3 => n2693, A4 => 
                           n2694, ZN => n2681);
   U2638 : AOI221_X1 port map( B1 => n662, B2 => n4996, C1 => n665, C2 => n5028
                           , A => n2695, ZN => n2694);
   U2639 : OAI22_X1 port map( A1 => n1815, A2 => n668, B1 => n1816, B2 => n671,
                           ZN => n2695);
   U2640 : AOI221_X1 port map( B1 => n674, B2 => n5284, C1 => n677, C2 => n5252
                           , A => n2696, ZN => n2693);
   U2641 : OAI22_X1 port map( A1 => n1818, A2 => n680, B1 => n1819, B2 => n683,
                           ZN => n2696);
   U2642 : AOI221_X1 port map( B1 => n686, B2 => n4548, C1 => n689, C2 => n4580
                           , A => n2697, ZN => n2692);
   U2643 : OAI22_X1 port map( A1 => n1821, A2 => n692, B1 => n1822, B2 => n695,
                           ZN => n2697);
   U2644 : AOI221_X1 port map( B1 => n698, B2 => n4612, C1 => n701, C2 => n4644
                           , A => n2698, ZN => n2691);
   U2645 : OAI22_X1 port map( A1 => n1824, A2 => n704, B1 => n1825, B2 => n707,
                           ZN => n2698);
   U2646 : NAND2_X1 port map( A1 => DATAIN(16), A2 => n264, ZN => n1797);
   U2647 : OAI21_X1 port map( B1 => n269, B2 => n2699, A => n711, ZN => n3015);
   U2648 : OAI221_X1 port map( B1 => n1827, B2 => n608, C1 => n274, C2 => n2700
                           , A => n2701, ZN => n3014);
   U2649 : OAI21_X1 port map( B1 => n2702, B2 => n2703, A => n611, ZN => n2701)
                           ;
   U2650 : NAND4_X1 port map( A1 => n2704, A2 => n2705, A3 => n2706, A4 => 
                           n2707, ZN => n2703);
   U2651 : AOI221_X1 port map( B1 => n614, B2 => n1046, C1 => n617, C2 => n1012
                           , A => n2708, ZN => n2707);
   U2652 : OAI22_X1 port map( A1 => n5059, A2 => n620, B1 => n5091, B2 => n623,
                           ZN => n2708);
   U2653 : AOI221_X1 port map( B1 => n626, B2 => n874, C1 => n629, C2 => n908, 
                           A => n2709, ZN => n2706);
   U2654 : OAI22_X1 port map( A1 => n5347, A2 => n632, B1 => n5315, B2 => n635,
                           ZN => n2709);
   U2655 : AOI221_X1 port map( B1 => n638, B2 => n1826, C1 => n641, C2 => n1295
                           , A => n2710, ZN => n2705);
   U2656 : OAI22_X1 port map( A1 => n4483, A2 => n644, B1 => n4515, B2 => n647,
                           ZN => n2710);
   U2657 : AOI221_X1 port map( B1 => n650, B2 => n1116, C1 => n653, C2 => n1082
                           , A => n2711, ZN => n2704);
   U2658 : OAI22_X1 port map( A1 => n4675, A2 => n656, B1 => n4707, B2 => n659,
                           ZN => n2711);
   U2659 : NAND4_X1 port map( A1 => n2712, A2 => n2713, A3 => n2714, A4 => 
                           n2715, ZN => n2702);
   U2660 : AOI221_X1 port map( B1 => n662, B2 => n4995, C1 => n665, C2 => n5027
                           , A => n2716, ZN => n2715);
   U2661 : OAI22_X1 port map( A1 => n1845, A2 => n668, B1 => n1846, B2 => n671,
                           ZN => n2716);
   U2662 : AOI221_X1 port map( B1 => n674, B2 => n5283, C1 => n677, C2 => n5251
                           , A => n2717, ZN => n2714);
   U2663 : OAI22_X1 port map( A1 => n1848, A2 => n680, B1 => n1849, B2 => n683,
                           ZN => n2717);
   U2664 : AOI221_X1 port map( B1 => n686, B2 => n4547, C1 => n689, C2 => n4579
                           , A => n2718, ZN => n2713);
   U2665 : OAI22_X1 port map( A1 => n1851, A2 => n692, B1 => n1852, B2 => n695,
                           ZN => n2718);
   U2666 : AOI221_X1 port map( B1 => n698, B2 => n4611, C1 => n701, C2 => n4643
                           , A => n2719, ZN => n2712);
   U2667 : OAI22_X1 port map( A1 => n1854, A2 => n704, B1 => n1855, B2 => n707,
                           ZN => n2719);
   U2668 : NAND2_X1 port map( A1 => DATAIN(15), A2 => n264, ZN => n1827);
   U2669 : OAI21_X1 port map( B1 => n270, B2 => n2720, A => n711, ZN => n3013);
   U2670 : OAI221_X1 port map( B1 => n1857, B2 => n608, C1 => n274, C2 => n2721
                           , A => n2722, ZN => n3012);
   U2671 : OAI21_X1 port map( B1 => n2723, B2 => n2724, A => n611, ZN => n2722)
                           ;
   U2672 : NAND4_X1 port map( A1 => n2725, A2 => n2726, A3 => n2855, A4 => 
                           n2856, ZN => n2724);
   U2673 : AOI221_X1 port map( B1 => n614, B2 => n1047, C1 => n617, C2 => n1013
                           , A => n2857, ZN => n2856);
   U2674 : OAI22_X1 port map( A1 => n5058, A2 => n620, B1 => n5090, B2 => n623,
                           ZN => n2857);
   U2675 : AOI221_X1 port map( B1 => n626, B2 => n875, C1 => n629, C2 => n909, 
                           A => n2858, ZN => n2855);
   U2676 : OAI22_X1 port map( A1 => n5346, A2 => n632, B1 => n5314, B2 => n635,
                           ZN => n2858);
   U2677 : AOI221_X1 port map( B1 => n638, B2 => n1856, C1 => n641, C2 => n1296
                           , A => n2859, ZN => n2726);
   U2678 : OAI22_X1 port map( A1 => n4482, A2 => n644, B1 => n4514, B2 => n647,
                           ZN => n2859);
   U2679 : AOI221_X1 port map( B1 => n650, B2 => n1117, C1 => n653, C2 => n1083
                           , A => n2860, ZN => n2725);
   U2680 : OAI22_X1 port map( A1 => n4674, A2 => n656, B1 => n4706, B2 => n659,
                           ZN => n2860);
   U2681 : NAND4_X1 port map( A1 => n2861, A2 => n2862, A3 => n2863, A4 => 
                           n2864, ZN => n2723);
   U2682 : AOI221_X1 port map( B1 => n662, B2 => n4994, C1 => n665, C2 => n5026
                           , A => n2865, ZN => n2864);
   U2683 : OAI22_X1 port map( A1 => n1875, A2 => n668, B1 => n1876, B2 => n671,
                           ZN => n2865);
   U2684 : AOI221_X1 port map( B1 => n674, B2 => n5282, C1 => n677, C2 => n5250
                           , A => n2866, ZN => n2863);
   U2685 : OAI22_X1 port map( A1 => n1878, A2 => n680, B1 => n1879, B2 => n683,
                           ZN => n2866);
   U2686 : AOI221_X1 port map( B1 => n686, B2 => n4546, C1 => n689, C2 => n4578
                           , A => n2867, ZN => n2862);
   U2687 : OAI22_X1 port map( A1 => n1881, A2 => n692, B1 => n1882, B2 => n695,
                           ZN => n2867);
   U2688 : AOI221_X1 port map( B1 => n698, B2 => n4610, C1 => n701, C2 => n4642
                           , A => n2868, ZN => n2861);
   U2689 : OAI22_X1 port map( A1 => n1884, A2 => n704, B1 => n1885, B2 => n707,
                           ZN => n2868);
   U2690 : NAND2_X1 port map( A1 => DATAIN(14), A2 => n264, ZN => n1857);
   U2691 : OAI21_X1 port map( B1 => n269, B2 => n2869, A => n711, ZN => n3011);
   U2692 : OAI221_X1 port map( B1 => n1887, B2 => n608, C1 => n275, C2 => n2870
                           , A => n2871, ZN => n3010);
   U2693 : OAI21_X1 port map( B1 => n2872, B2 => n2873, A => n611, ZN => n2871)
                           ;
   U2694 : NAND4_X1 port map( A1 => n2874, A2 => n2875, A3 => n2876, A4 => 
                           n2877, ZN => n2873);
   U2695 : AOI221_X1 port map( B1 => n614, B2 => n1048, C1 => n617, C2 => n1014
                           , A => n2878, ZN => n2877);
   U2696 : OAI22_X1 port map( A1 => n5057, A2 => n620, B1 => n5089, B2 => n623,
                           ZN => n2878);
   U2697 : AOI221_X1 port map( B1 => n626, B2 => n876, C1 => n629, C2 => n910, 
                           A => n2879, ZN => n2876);
   U2698 : OAI22_X1 port map( A1 => n5345, A2 => n632, B1 => n5313, B2 => n635,
                           ZN => n2879);
   U2699 : AOI221_X1 port map( B1 => n638, B2 => n1886, C1 => n641, C2 => n1297
                           , A => n2880, ZN => n2875);
   U2700 : OAI22_X1 port map( A1 => n4481, A2 => n644, B1 => n4513, B2 => n647,
                           ZN => n2880);
   U2701 : AOI221_X1 port map( B1 => n650, B2 => n1118, C1 => n653, C2 => n1084
                           , A => n2881, ZN => n2874);
   U2702 : OAI22_X1 port map( A1 => n4673, A2 => n656, B1 => n4705, B2 => n659,
                           ZN => n2881);
   U2703 : NAND4_X1 port map( A1 => n2882, A2 => n2883, A3 => n2884, A4 => 
                           n2885, ZN => n2872);
   U2704 : AOI221_X1 port map( B1 => n662, B2 => n4993, C1 => n665, C2 => n5025
                           , A => n2886, ZN => n2885);
   U2705 : OAI22_X1 port map( A1 => n1905, A2 => n668, B1 => n1906, B2 => n671,
                           ZN => n2886);
   U2706 : AOI221_X1 port map( B1 => n674, B2 => n5281, C1 => n677, C2 => n5249
                           , A => n2887, ZN => n2884);
   U2707 : OAI22_X1 port map( A1 => n1908, A2 => n680, B1 => n1909, B2 => n683,
                           ZN => n2887);
   U2708 : AOI221_X1 port map( B1 => n686, B2 => n4545, C1 => n689, C2 => n4577
                           , A => n2888, ZN => n2883);
   U2709 : OAI22_X1 port map( A1 => n1911, A2 => n692, B1 => n1912, B2 => n695,
                           ZN => n2888);
   U2710 : AOI221_X1 port map( B1 => n698, B2 => n4609, C1 => n701, C2 => n4641
                           , A => n2889, ZN => n2882);
   U2711 : OAI22_X1 port map( A1 => n1914, A2 => n704, B1 => n1915, B2 => n707,
                           ZN => n2889);
   U2712 : NAND2_X1 port map( A1 => DATAIN(13), A2 => n263, ZN => n1887);
   U2713 : OAI21_X1 port map( B1 => n270, B2 => n2890, A => n711, ZN => n3009);
   U2714 : OAI221_X1 port map( B1 => n1917, B2 => n608, C1 => n274, C2 => n2891
                           , A => n2892, ZN => n3008);
   U2715 : OAI21_X1 port map( B1 => n2893, B2 => n2894, A => n611, ZN => n2892)
                           ;
   U2716 : NAND4_X1 port map( A1 => n2895, A2 => n2896, A3 => n2897, A4 => 
                           n2898, ZN => n2894);
   U2717 : AOI221_X1 port map( B1 => n614, B2 => n1049, C1 => n617, C2 => n1015
                           , A => n2899, ZN => n2898);
   U2718 : OAI22_X1 port map( A1 => n5056, A2 => n620, B1 => n5088, B2 => n623,
                           ZN => n2899);
   U2719 : AOI221_X1 port map( B1 => n626, B2 => n877, C1 => n629, C2 => n911, 
                           A => n2900, ZN => n2897);
   U2720 : OAI22_X1 port map( A1 => n5344, A2 => n632, B1 => n5312, B2 => n635,
                           ZN => n2900);
   U2721 : AOI221_X1 port map( B1 => n638, B2 => n1916, C1 => n641, C2 => n1298
                           , A => n2901, ZN => n2896);
   U2722 : OAI22_X1 port map( A1 => n4480, A2 => n644, B1 => n4512, B2 => n647,
                           ZN => n2901);
   U2723 : AOI221_X1 port map( B1 => n650, B2 => n1119, C1 => n653, C2 => n1085
                           , A => n2902, ZN => n2895);
   U2724 : OAI22_X1 port map( A1 => n4672, A2 => n656, B1 => n4704, B2 => n659,
                           ZN => n2902);
   U2725 : NAND4_X1 port map( A1 => n2903, A2 => n2904, A3 => n2905, A4 => 
                           n2906, ZN => n2893);
   U2726 : AOI221_X1 port map( B1 => n662, B2 => n4992, C1 => n665, C2 => n5024
                           , A => n2907, ZN => n2906);
   U2727 : OAI22_X1 port map( A1 => n1935, A2 => n668, B1 => n1936, B2 => n671,
                           ZN => n2907);
   U2728 : AOI221_X1 port map( B1 => n674, B2 => n5280, C1 => n677, C2 => n5248
                           , A => n2908, ZN => n2905);
   U2729 : OAI22_X1 port map( A1 => n1938, A2 => n680, B1 => n1939, B2 => n683,
                           ZN => n2908);
   U2730 : AOI221_X1 port map( B1 => n686, B2 => n4544, C1 => n689, C2 => n4576
                           , A => n2909, ZN => n2904);
   U2731 : OAI22_X1 port map( A1 => n1941, A2 => n692, B1 => n1942, B2 => n695,
                           ZN => n2909);
   U2732 : AOI221_X1 port map( B1 => n698, B2 => n4608, C1 => n701, C2 => n4640
                           , A => n2910, ZN => n2903);
   U2733 : OAI22_X1 port map( A1 => n1944, A2 => n704, B1 => n1945, B2 => n707,
                           ZN => n2910);
   U2734 : NAND2_X1 port map( A1 => DATAIN(12), A2 => n263, ZN => n1917);
   U2735 : OAI21_X1 port map( B1 => n269, B2 => n2911, A => n711, ZN => n3007);
   U2736 : OAI221_X1 port map( B1 => n1947, B2 => n608, C1 => n274, C2 => n2912
                           , A => n2913, ZN => n3006);
   U2737 : OAI21_X1 port map( B1 => n2914, B2 => n2915, A => n610, ZN => n2913)
                           ;
   U2738 : NAND4_X1 port map( A1 => n2916, A2 => n2917, A3 => n2918, A4 => 
                           n2919, ZN => n2915);
   U2739 : AOI221_X1 port map( B1 => n613, B2 => n1050, C1 => n616, C2 => n1016
                           , A => n2920, ZN => n2919);
   U2740 : OAI22_X1 port map( A1 => n5055, A2 => n619, B1 => n5087, B2 => n622,
                           ZN => n2920);
   U2741 : AOI221_X1 port map( B1 => n625, B2 => n878, C1 => n628, C2 => n912, 
                           A => n2921, ZN => n2918);
   U2742 : OAI22_X1 port map( A1 => n5343, A2 => n631, B1 => n5311, B2 => n634,
                           ZN => n2921);
   U2743 : AOI221_X1 port map( B1 => n637, B2 => n1946, C1 => n640, C2 => n1299
                           , A => n2922, ZN => n2917);
   U2744 : OAI22_X1 port map( A1 => n4479, A2 => n643, B1 => n4511, B2 => n646,
                           ZN => n2922);
   U2745 : AOI221_X1 port map( B1 => n649, B2 => n1120, C1 => n652, C2 => n1086
                           , A => n2923, ZN => n2916);
   U2746 : OAI22_X1 port map( A1 => n4671, A2 => n655, B1 => n4703, B2 => n658,
                           ZN => n2923);
   U2747 : NAND4_X1 port map( A1 => n2924, A2 => n2925, A3 => n2926, A4 => 
                           n2927, ZN => n2914);
   U2748 : AOI221_X1 port map( B1 => n661, B2 => n4991, C1 => n664, C2 => n5023
                           , A => n2928, ZN => n2927);
   U2749 : OAI22_X1 port map( A1 => n1965, A2 => n667, B1 => n1966, B2 => n670,
                           ZN => n2928);
   U2750 : AOI221_X1 port map( B1 => n673, B2 => n5279, C1 => n676, C2 => n5247
                           , A => n2929, ZN => n2926);
   U2751 : OAI22_X1 port map( A1 => n1968, A2 => n679, B1 => n1969, B2 => n682,
                           ZN => n2929);
   U2752 : AOI221_X1 port map( B1 => n685, B2 => n4543, C1 => n688, C2 => n4575
                           , A => n2930, ZN => n2925);
   U2753 : OAI22_X1 port map( A1 => n1971, A2 => n691, B1 => n1972, B2 => n694,
                           ZN => n2930);
   U2754 : AOI221_X1 port map( B1 => n697, B2 => n4607, C1 => n700, C2 => n4639
                           , A => n2931, ZN => n2924);
   U2755 : OAI22_X1 port map( A1 => n1974, A2 => n703, B1 => n1975, B2 => n706,
                           ZN => n2931);
   U2756 : NAND2_X1 port map( A1 => DATAIN(11), A2 => n263, ZN => n1947);
   U2757 : OAI21_X1 port map( B1 => n270, B2 => n2932, A => n710, ZN => n3005);
   U2758 : OAI221_X1 port map( B1 => n1977, B2 => n608, C1 => n274, C2 => n2933
                           , A => n2934, ZN => n3004);
   U2759 : OAI21_X1 port map( B1 => n2935, B2 => n2936, A => n610, ZN => n2934)
                           ;
   U2760 : NAND4_X1 port map( A1 => n2937, A2 => n2938, A3 => n2939, A4 => 
                           n2940, ZN => n2936);
   U2761 : AOI221_X1 port map( B1 => n613, B2 => n1051, C1 => n616, C2 => n1017
                           , A => n2941, ZN => n2940);
   U2762 : OAI22_X1 port map( A1 => n5054, A2 => n619, B1 => n5086, B2 => n622,
                           ZN => n2941);
   U2763 : AOI221_X1 port map( B1 => n625, B2 => n879, C1 => n628, C2 => n913, 
                           A => n2942, ZN => n2939);
   U2764 : OAI22_X1 port map( A1 => n5342, A2 => n631, B1 => n5310, B2 => n634,
                           ZN => n2942);
   U2765 : AOI221_X1 port map( B1 => n637, B2 => n1976, C1 => n640, C2 => n1300
                           , A => n2943, ZN => n2938);
   U2766 : OAI22_X1 port map( A1 => n4478, A2 => n643, B1 => n4510, B2 => n646,
                           ZN => n2943);
   U2767 : AOI221_X1 port map( B1 => n649, B2 => n1121, C1 => n652, C2 => n1087
                           , A => n2944, ZN => n2937);
   U2768 : OAI22_X1 port map( A1 => n4670, A2 => n655, B1 => n4702, B2 => n658,
                           ZN => n2944);
   U2769 : NAND4_X1 port map( A1 => n2945, A2 => n2946, A3 => n2947, A4 => 
                           n2948, ZN => n2935);
   U2770 : AOI221_X1 port map( B1 => n661, B2 => n4990, C1 => n664, C2 => n5022
                           , A => n2949, ZN => n2948);
   U2771 : OAI22_X1 port map( A1 => n1995, A2 => n667, B1 => n1996, B2 => n670,
                           ZN => n2949);
   U2772 : AOI221_X1 port map( B1 => n673, B2 => n5278, C1 => n676, C2 => n5246
                           , A => n2950, ZN => n2947);
   U2773 : OAI22_X1 port map( A1 => n1998, A2 => n679, B1 => n1999, B2 => n682,
                           ZN => n2950);
   U2774 : AOI221_X1 port map( B1 => n685, B2 => n4542, C1 => n688, C2 => n4574
                           , A => n2951, ZN => n2946);
   U2775 : OAI22_X1 port map( A1 => n2001, A2 => n691, B1 => n2002, B2 => n694,
                           ZN => n2951);
   U2776 : AOI221_X1 port map( B1 => n697, B2 => n4606, C1 => n700, C2 => n4638
                           , A => n2952, ZN => n2945);
   U2777 : OAI22_X1 port map( A1 => n2004, A2 => n703, B1 => n2005, B2 => n706,
                           ZN => n2952);
   U2778 : NAND2_X1 port map( A1 => DATAIN(10), A2 => n263, ZN => n1977);
   U2779 : OAI21_X1 port map( B1 => n269, B2 => n2953, A => n710, ZN => n3003);
   U2780 : OAI221_X1 port map( B1 => n2007, B2 => n608, C1 => n274, C2 => n2954
                           , A => n2955, ZN => n3002);
   U2781 : OAI21_X1 port map( B1 => n2956, B2 => n2957, A => n610, ZN => n2955)
                           ;
   U2782 : NAND4_X1 port map( A1 => n2958, A2 => n2959, A3 => n2960, A4 => 
                           n2961, ZN => n2957);
   U2783 : AOI221_X1 port map( B1 => n613, B2 => n1052, C1 => n616, C2 => n1018
                           , A => n2962, ZN => n2961);
   U2784 : OAI22_X1 port map( A1 => n5053, A2 => n619, B1 => n5085, B2 => n622,
                           ZN => n2962);
   U2785 : AOI221_X1 port map( B1 => n625, B2 => n880, C1 => n628, C2 => n914, 
                           A => n2963, ZN => n2960);
   U2786 : OAI22_X1 port map( A1 => n5341, A2 => n631, B1 => n5309, B2 => n634,
                           ZN => n2963);
   U2787 : AOI221_X1 port map( B1 => n637, B2 => n2006, C1 => n640, C2 => n1301
                           , A => n2964, ZN => n2959);
   U2788 : OAI22_X1 port map( A1 => n4477, A2 => n643, B1 => n4509, B2 => n646,
                           ZN => n2964);
   U2789 : AOI221_X1 port map( B1 => n649, B2 => n1122, C1 => n652, C2 => n1088
                           , A => n2965, ZN => n2958);
   U2790 : OAI22_X1 port map( A1 => n4669, A2 => n655, B1 => n4701, B2 => n658,
                           ZN => n2965);
   U2791 : NAND4_X1 port map( A1 => n2966, A2 => n2967, A3 => n2968, A4 => 
                           n2969, ZN => n2956);
   U2792 : AOI221_X1 port map( B1 => n661, B2 => n4989, C1 => n664, C2 => n5021
                           , A => n2970, ZN => n2969);
   U2793 : OAI22_X1 port map( A1 => n2025, A2 => n667, B1 => n2026, B2 => n670,
                           ZN => n2970);
   U2794 : AOI221_X1 port map( B1 => n673, B2 => n5277, C1 => n676, C2 => n5245
                           , A => n2971, ZN => n2968);
   U2795 : OAI22_X1 port map( A1 => n2028, A2 => n679, B1 => n2029, B2 => n682,
                           ZN => n2971);
   U2796 : AOI221_X1 port map( B1 => n685, B2 => n4541, C1 => n688, C2 => n4573
                           , A => n2972, ZN => n2967);
   U2797 : OAI22_X1 port map( A1 => n2031, A2 => n691, B1 => n2032, B2 => n694,
                           ZN => n2972);
   U2798 : AOI221_X1 port map( B1 => n697, B2 => n4605, C1 => n700, C2 => n4637
                           , A => n2973, ZN => n2966);
   U2799 : OAI22_X1 port map( A1 => n2034, A2 => n703, B1 => n2035, B2 => n706,
                           ZN => n2973);
   U2800 : NAND2_X1 port map( A1 => DATAIN(9), A2 => n263, ZN => n2007);
   U2801 : OAI21_X1 port map( B1 => n268, B2 => n2974, A => n710, ZN => n3001);
   U2802 : OAI221_X1 port map( B1 => n2037, B2 => n608, C1 => n275, C2 => n2975
                           , A => n2976, ZN => n3000);
   U2803 : OAI21_X1 port map( B1 => n2977, B2 => n2978, A => n610, ZN => n2976)
                           ;
   U2804 : NAND4_X1 port map( A1 => n2979, A2 => n2980, A3 => n2981, A4 => 
                           n2982, ZN => n2978);
   U2805 : AOI221_X1 port map( B1 => n613, B2 => n1053, C1 => n616, C2 => n1019
                           , A => n4135, ZN => n2982);
   U2806 : OAI22_X1 port map( A1 => n5052, A2 => n619, B1 => n5084, B2 => n622,
                           ZN => n4135);
   U2807 : AOI221_X1 port map( B1 => n625, B2 => n881, C1 => n628, C2 => n915, 
                           A => n4136, ZN => n2981);
   U2808 : OAI22_X1 port map( A1 => n5340, A2 => n631, B1 => n5308, B2 => n634,
                           ZN => n4136);
   U2809 : AOI221_X1 port map( B1 => n637, B2 => n2036, C1 => n640, C2 => n1302
                           , A => n4137, ZN => n2980);
   U2810 : OAI22_X1 port map( A1 => n4476, A2 => n643, B1 => n4508, B2 => n646,
                           ZN => n4137);
   U2811 : AOI221_X1 port map( B1 => n649, B2 => n1123, C1 => n652, C2 => n1089
                           , A => n4138, ZN => n2979);
   U2812 : OAI22_X1 port map( A1 => n4668, A2 => n655, B1 => n4700, B2 => n658,
                           ZN => n4138);
   U2813 : NAND4_X1 port map( A1 => n4139, A2 => n4140, A3 => n4141, A4 => 
                           n4142, ZN => n2977);
   U2814 : AOI221_X1 port map( B1 => n661, B2 => n4988, C1 => n664, C2 => n5020
                           , A => n4143, ZN => n4142);
   U2815 : OAI22_X1 port map( A1 => n2055, A2 => n667, B1 => n2056, B2 => n670,
                           ZN => n4143);
   U2816 : AOI221_X1 port map( B1 => n673, B2 => n5276, C1 => n676, C2 => n5244
                           , A => n4144, ZN => n4141);
   U2817 : OAI22_X1 port map( A1 => n2058, A2 => n679, B1 => n2059, B2 => n682,
                           ZN => n4144);
   U2818 : AOI221_X1 port map( B1 => n685, B2 => n4540, C1 => n688, C2 => n4572
                           , A => n4145, ZN => n4140);
   U2819 : OAI22_X1 port map( A1 => n2061, A2 => n691, B1 => n2062, B2 => n694,
                           ZN => n4145);
   U2820 : AOI221_X1 port map( B1 => n697, B2 => n4604, C1 => n700, C2 => n4636
                           , A => n4146, ZN => n4139);
   U2821 : OAI22_X1 port map( A1 => n2064, A2 => n703, B1 => n2065, B2 => n706,
                           ZN => n4146);
   U2822 : NAND2_X1 port map( A1 => DATAIN(8), A2 => n263, ZN => n2037);
   U2823 : OAI21_X1 port map( B1 => n269, B2 => n4147, A => n710, ZN => n2999);
   U2824 : OAI221_X1 port map( B1 => n2067, B2 => n609, C1 => n275, C2 => n4148
                           , A => n4149, ZN => n2998);
   U2825 : OAI21_X1 port map( B1 => n4150, B2 => n4151, A => n610, ZN => n4149)
                           ;
   U2826 : NAND4_X1 port map( A1 => n4152, A2 => n4153, A3 => n4154, A4 => 
                           n4155, ZN => n4151);
   U2827 : AOI221_X1 port map( B1 => n613, B2 => n1054, C1 => n616, C2 => n1020
                           , A => n4156, ZN => n4155);
   U2828 : OAI22_X1 port map( A1 => n5051, A2 => n619, B1 => n5083, B2 => n622,
                           ZN => n4156);
   U2829 : AOI221_X1 port map( B1 => n625, B2 => n882, C1 => n628, C2 => n916, 
                           A => n4157, ZN => n4154);
   U2830 : OAI22_X1 port map( A1 => n5339, A2 => n631, B1 => n5307, B2 => n634,
                           ZN => n4157);
   U2831 : AOI221_X1 port map( B1 => n637, B2 => n2066, C1 => n640, C2 => n1303
                           , A => n4158, ZN => n4153);
   U2832 : OAI22_X1 port map( A1 => n4475, A2 => n643, B1 => n4507, B2 => n646,
                           ZN => n4158);
   U2833 : AOI221_X1 port map( B1 => n649, B2 => n1124, C1 => n652, C2 => n1090
                           , A => n4159, ZN => n4152);
   U2834 : OAI22_X1 port map( A1 => n4667, A2 => n655, B1 => n4699, B2 => n658,
                           ZN => n4159);
   U2835 : NAND4_X1 port map( A1 => n4160, A2 => n4161, A3 => n4162, A4 => 
                           n4163, ZN => n4150);
   U2836 : AOI221_X1 port map( B1 => n661, B2 => n4987, C1 => n664, C2 => n5019
                           , A => n4164, ZN => n4163);
   U2837 : OAI22_X1 port map( A1 => n2085, A2 => n667, B1 => n2086, B2 => n670,
                           ZN => n4164);
   U2838 : AOI221_X1 port map( B1 => n673, B2 => n5275, C1 => n676, C2 => n5243
                           , A => n4165, ZN => n4162);
   U2839 : OAI22_X1 port map( A1 => n2088, A2 => n679, B1 => n2089, B2 => n682,
                           ZN => n4165);
   U2840 : AOI221_X1 port map( B1 => n685, B2 => n4539, C1 => n688, C2 => n4571
                           , A => n4166, ZN => n4161);
   U2841 : OAI22_X1 port map( A1 => n2091, A2 => n691, B1 => n2092, B2 => n694,
                           ZN => n4166);
   U2842 : AOI221_X1 port map( B1 => n697, B2 => n4603, C1 => n700, C2 => n4635
                           , A => n4167, ZN => n4160);
   U2843 : OAI22_X1 port map( A1 => n2094, A2 => n703, B1 => n2095, B2 => n706,
                           ZN => n4167);
   U2844 : NAND2_X1 port map( A1 => DATAIN(7), A2 => n263, ZN => n2067);
   U2845 : OAI21_X1 port map( B1 => n270, B2 => n4168, A => n710, ZN => n2997);
   U2846 : OAI221_X1 port map( B1 => n2097, B2 => n609, C1 => n275, C2 => n4169
                           , A => n4170, ZN => n2996);
   U2847 : OAI21_X1 port map( B1 => n4171, B2 => n4172, A => n610, ZN => n4170)
                           ;
   U2848 : NAND4_X1 port map( A1 => n4173, A2 => n4174, A3 => n4175, A4 => 
                           n4176, ZN => n4172);
   U2849 : AOI221_X1 port map( B1 => n613, B2 => n1055, C1 => n616, C2 => n1021
                           , A => n4177, ZN => n4176);
   U2850 : OAI22_X1 port map( A1 => n5050, A2 => n619, B1 => n5082, B2 => n622,
                           ZN => n4177);
   U2851 : AOI221_X1 port map( B1 => n625, B2 => n883, C1 => n628, C2 => n917, 
                           A => n4178, ZN => n4175);
   U2852 : OAI22_X1 port map( A1 => n5338, A2 => n631, B1 => n5306, B2 => n634,
                           ZN => n4178);
   U2853 : AOI221_X1 port map( B1 => n637, B2 => n2096, C1 => n640, C2 => n1304
                           , A => n4179, ZN => n4174);
   U2854 : OAI22_X1 port map( A1 => n4474, A2 => n643, B1 => n4506, B2 => n646,
                           ZN => n4179);
   U2855 : AOI221_X1 port map( B1 => n649, B2 => n1125, C1 => n652, C2 => n1091
                           , A => n4180, ZN => n4173);
   U2856 : OAI22_X1 port map( A1 => n4666, A2 => n655, B1 => n4698, B2 => n658,
                           ZN => n4180);
   U2857 : NAND4_X1 port map( A1 => n4181, A2 => n4182, A3 => n4183, A4 => 
                           n4184, ZN => n4171);
   U2858 : AOI221_X1 port map( B1 => n661, B2 => n4986, C1 => n664, C2 => n5018
                           , A => n4185, ZN => n4184);
   U2859 : OAI22_X1 port map( A1 => n2115, A2 => n667, B1 => n2116, B2 => n670,
                           ZN => n4185);
   U2860 : AOI221_X1 port map( B1 => n673, B2 => n5274, C1 => n676, C2 => n5242
                           , A => n4186, ZN => n4183);
   U2861 : OAI22_X1 port map( A1 => n2118, A2 => n679, B1 => n2119, B2 => n682,
                           ZN => n4186);
   U2862 : AOI221_X1 port map( B1 => n685, B2 => n4538, C1 => n688, C2 => n4570
                           , A => n4187, ZN => n4182);
   U2863 : OAI22_X1 port map( A1 => n2121, A2 => n691, B1 => n2122, B2 => n694,
                           ZN => n4187);
   U2864 : AOI221_X1 port map( B1 => n697, B2 => n4602, C1 => n700, C2 => n4634
                           , A => n4188, ZN => n4181);
   U2865 : OAI22_X1 port map( A1 => n2124, A2 => n703, B1 => n2125, B2 => n706,
                           ZN => n4188);
   U2866 : NAND2_X1 port map( A1 => DATAIN(6), A2 => n263, ZN => n2097);
   U2867 : OAI21_X1 port map( B1 => n269, B2 => n4189, A => n710, ZN => n2995);
   U2868 : OAI221_X1 port map( B1 => n2127, B2 => n609, C1 => n275, C2 => n4190
                           , A => n4191, ZN => n2994);
   U2869 : OAI21_X1 port map( B1 => n4192, B2 => n4193, A => n610, ZN => n4191)
                           ;
   U2870 : NAND4_X1 port map( A1 => n4194, A2 => n4195, A3 => n4196, A4 => 
                           n4197, ZN => n4193);
   U2871 : AOI221_X1 port map( B1 => n613, B2 => n1056, C1 => n616, C2 => n1022
                           , A => n4198, ZN => n4197);
   U2872 : OAI22_X1 port map( A1 => n5049, A2 => n619, B1 => n5081, B2 => n622,
                           ZN => n4198);
   U2873 : AOI221_X1 port map( B1 => n625, B2 => n884, C1 => n628, C2 => n918, 
                           A => n4199, ZN => n4196);
   U2874 : OAI22_X1 port map( A1 => n5337, A2 => n631, B1 => n5305, B2 => n634,
                           ZN => n4199);
   U2875 : AOI221_X1 port map( B1 => n637, B2 => n2126, C1 => n640, C2 => n1305
                           , A => n4200, ZN => n4195);
   U2876 : OAI22_X1 port map( A1 => n4473, A2 => n643, B1 => n4505, B2 => n646,
                           ZN => n4200);
   U2877 : AOI221_X1 port map( B1 => n649, B2 => n1126, C1 => n652, C2 => n1092
                           , A => n4201, ZN => n4194);
   U2878 : OAI22_X1 port map( A1 => n4665, A2 => n655, B1 => n4697, B2 => n658,
                           ZN => n4201);
   U2879 : NAND4_X1 port map( A1 => n4202, A2 => n4203, A3 => n4204, A4 => 
                           n4205, ZN => n4192);
   U2880 : AOI221_X1 port map( B1 => n661, B2 => n4985, C1 => n664, C2 => n5017
                           , A => n4206, ZN => n4205);
   U2881 : OAI22_X1 port map( A1 => n2145, A2 => n667, B1 => n2146, B2 => n670,
                           ZN => n4206);
   U2882 : AOI221_X1 port map( B1 => n673, B2 => n5273, C1 => n676, C2 => n5241
                           , A => n4207, ZN => n4204);
   U2883 : OAI22_X1 port map( A1 => n2148, A2 => n679, B1 => n2149, B2 => n682,
                           ZN => n4207);
   U2884 : AOI221_X1 port map( B1 => n685, B2 => n4537, C1 => n688, C2 => n4569
                           , A => n4208, ZN => n4203);
   U2885 : OAI22_X1 port map( A1 => n2151, A2 => n691, B1 => n2152, B2 => n694,
                           ZN => n4208);
   U2886 : AOI221_X1 port map( B1 => n697, B2 => n4601, C1 => n700, C2 => n4633
                           , A => n4209, ZN => n4202);
   U2887 : OAI22_X1 port map( A1 => n2154, A2 => n703, B1 => n2155, B2 => n706,
                           ZN => n4209);
   U2888 : NAND2_X1 port map( A1 => DATAIN(5), A2 => n263, ZN => n2127);
   U2889 : OAI21_X1 port map( B1 => n270, B2 => n4210, A => n710, ZN => n2993);
   U2890 : OAI221_X1 port map( B1 => n2157, B2 => n609, C1 => n275, C2 => n4211
                           , A => n4212, ZN => n2992);
   U2891 : OAI21_X1 port map( B1 => n4213, B2 => n4214, A => n610, ZN => n4212)
                           ;
   U2892 : NAND4_X1 port map( A1 => n4215, A2 => n4216, A3 => n4217, A4 => 
                           n4218, ZN => n4214);
   U2893 : AOI221_X1 port map( B1 => n613, B2 => n1057, C1 => n616, C2 => n1023
                           , A => n4219, ZN => n4218);
   U2894 : OAI22_X1 port map( A1 => n5048, A2 => n619, B1 => n5080, B2 => n622,
                           ZN => n4219);
   U2895 : AOI221_X1 port map( B1 => n625, B2 => n885, C1 => n628, C2 => n919, 
                           A => n4220, ZN => n4217);
   U2896 : OAI22_X1 port map( A1 => n5336, A2 => n631, B1 => n5304, B2 => n634,
                           ZN => n4220);
   U2897 : AOI221_X1 port map( B1 => n637, B2 => n2156, C1 => n640, C2 => n1306
                           , A => n4221, ZN => n4216);
   U2898 : OAI22_X1 port map( A1 => n4472, A2 => n643, B1 => n4504, B2 => n646,
                           ZN => n4221);
   U2899 : AOI221_X1 port map( B1 => n649, B2 => n1127, C1 => n652, C2 => n1093
                           , A => n4222, ZN => n4215);
   U2900 : OAI22_X1 port map( A1 => n4664, A2 => n655, B1 => n4696, B2 => n658,
                           ZN => n4222);
   U2901 : NAND4_X1 port map( A1 => n4223, A2 => n4224, A3 => n4225, A4 => 
                           n4226, ZN => n4213);
   U2902 : AOI221_X1 port map( B1 => n661, B2 => n4984, C1 => n664, C2 => n5016
                           , A => n4227, ZN => n4226);
   U2903 : OAI22_X1 port map( A1 => n2175, A2 => n667, B1 => n2176, B2 => n670,
                           ZN => n4227);
   U2904 : AOI221_X1 port map( B1 => n673, B2 => n5272, C1 => n676, C2 => n5240
                           , A => n4228, ZN => n4225);
   U2905 : OAI22_X1 port map( A1 => n2178, A2 => n679, B1 => n2179, B2 => n682,
                           ZN => n4228);
   U2906 : AOI221_X1 port map( B1 => n685, B2 => n4536, C1 => n688, C2 => n4568
                           , A => n4229, ZN => n4224);
   U2907 : OAI22_X1 port map( A1 => n2181, A2 => n691, B1 => n2182, B2 => n694,
                           ZN => n4229);
   U2908 : AOI221_X1 port map( B1 => n697, B2 => n4600, C1 => n700, C2 => n4632
                           , A => n4230, ZN => n4223);
   U2909 : OAI22_X1 port map( A1 => n2184, A2 => n703, B1 => n2185, B2 => n706,
                           ZN => n4230);
   U2910 : NAND2_X1 port map( A1 => DATAIN(4), A2 => n263, ZN => n2157);
   U2911 : OAI21_X1 port map( B1 => n269, B2 => n4231, A => n710, ZN => n2991);
   U2912 : OAI221_X1 port map( B1 => n2187, B2 => n609, C1 => n275, C2 => n4232
                           , A => n4233, ZN => n2990);
   U2913 : OAI21_X1 port map( B1 => n4234, B2 => n4235, A => n610, ZN => n4233)
                           ;
   U2914 : NAND4_X1 port map( A1 => n4236, A2 => n4237, A3 => n4238, A4 => 
                           n4239, ZN => n4235);
   U2915 : AOI221_X1 port map( B1 => n613, B2 => n1058, C1 => n616, C2 => n1024
                           , A => n4240, ZN => n4239);
   U2916 : OAI22_X1 port map( A1 => n5047, A2 => n619, B1 => n5079, B2 => n622,
                           ZN => n4240);
   U2917 : AOI221_X1 port map( B1 => n625, B2 => n886, C1 => n628, C2 => n920, 
                           A => n4241, ZN => n4238);
   U2918 : OAI22_X1 port map( A1 => n5335, A2 => n631, B1 => n5303, B2 => n634,
                           ZN => n4241);
   U2919 : AOI221_X1 port map( B1 => n637, B2 => n2186, C1 => n640, C2 => n1307
                           , A => n4242, ZN => n4237);
   U2920 : OAI22_X1 port map( A1 => n4471, A2 => n643, B1 => n4503, B2 => n646,
                           ZN => n4242);
   U2921 : AOI221_X1 port map( B1 => n649, B2 => n1128, C1 => n652, C2 => n1094
                           , A => n4243, ZN => n4236);
   U2922 : OAI22_X1 port map( A1 => n4663, A2 => n655, B1 => n4695, B2 => n658,
                           ZN => n4243);
   U2923 : NAND4_X1 port map( A1 => n4244, A2 => n4245, A3 => n4246, A4 => 
                           n4247, ZN => n4234);
   U2924 : AOI221_X1 port map( B1 => n661, B2 => n4983, C1 => n664, C2 => n5015
                           , A => n4248, ZN => n4247);
   U2925 : OAI22_X1 port map( A1 => n2205, A2 => n667, B1 => n2206, B2 => n670,
                           ZN => n4248);
   U2926 : AOI221_X1 port map( B1 => n673, B2 => n5271, C1 => n676, C2 => n5239
                           , A => n4249, ZN => n4246);
   U2927 : OAI22_X1 port map( A1 => n2208, A2 => n679, B1 => n2209, B2 => n682,
                           ZN => n4249);
   U2928 : AOI221_X1 port map( B1 => n685, B2 => n4535, C1 => n688, C2 => n4567
                           , A => n4250, ZN => n4245);
   U2929 : OAI22_X1 port map( A1 => n2211, A2 => n691, B1 => n2212, B2 => n694,
                           ZN => n4250);
   U2930 : AOI221_X1 port map( B1 => n697, B2 => n4599, C1 => n700, C2 => n4631
                           , A => n4251, ZN => n4244);
   U2931 : OAI22_X1 port map( A1 => n2214, A2 => n703, B1 => n2215, B2 => n706,
                           ZN => n4251);
   U2932 : NAND2_X1 port map( A1 => DATAIN(3), A2 => n263, ZN => n2187);
   U2933 : OAI21_X1 port map( B1 => n270, B2 => n4252, A => n710, ZN => n2989);
   U2934 : OAI221_X1 port map( B1 => n2217, B2 => n609, C1 => n275, C2 => n4253
                           , A => n4254, ZN => n2988);
   U2935 : OAI21_X1 port map( B1 => n4255, B2 => n4256, A => n610, ZN => n4254)
                           ;
   U2936 : NAND4_X1 port map( A1 => n4257, A2 => n4258, A3 => n4259, A4 => 
                           n4260, ZN => n4256);
   U2937 : AOI221_X1 port map( B1 => n613, B2 => n1059, C1 => n616, C2 => n1025
                           , A => n4261, ZN => n4260);
   U2938 : OAI22_X1 port map( A1 => n5046, A2 => n619, B1 => n5078, B2 => n622,
                           ZN => n4261);
   U2939 : AOI221_X1 port map( B1 => n625, B2 => n887, C1 => n628, C2 => n921, 
                           A => n4262, ZN => n4259);
   U2940 : OAI22_X1 port map( A1 => n5334, A2 => n631, B1 => n5302, B2 => n634,
                           ZN => n4262);
   U2941 : AOI221_X1 port map( B1 => n637, B2 => n2216, C1 => n640, C2 => n1308
                           , A => n4263, ZN => n4258);
   U2942 : OAI22_X1 port map( A1 => n4470, A2 => n643, B1 => n4502, B2 => n646,
                           ZN => n4263);
   U2943 : AOI221_X1 port map( B1 => n649, B2 => n1129, C1 => n652, C2 => n1095
                           , A => n4264, ZN => n4257);
   U2944 : OAI22_X1 port map( A1 => n4662, A2 => n655, B1 => n4694, B2 => n658,
                           ZN => n4264);
   U2945 : NAND4_X1 port map( A1 => n4265, A2 => n4266, A3 => n4267, A4 => 
                           n4268, ZN => n4255);
   U2946 : AOI221_X1 port map( B1 => n661, B2 => n4982, C1 => n664, C2 => n5014
                           , A => n4269, ZN => n4268);
   U2947 : OAI22_X1 port map( A1 => n2235, A2 => n667, B1 => n2236, B2 => n670,
                           ZN => n4269);
   U2948 : AOI221_X1 port map( B1 => n673, B2 => n5270, C1 => n676, C2 => n5238
                           , A => n4270, ZN => n4267);
   U2949 : OAI22_X1 port map( A1 => n2238, A2 => n679, B1 => n2239, B2 => n682,
                           ZN => n4270);
   U2950 : AOI221_X1 port map( B1 => n685, B2 => n4534, C1 => n688, C2 => n4566
                           , A => n4271, ZN => n4266);
   U2951 : OAI22_X1 port map( A1 => n2241, A2 => n691, B1 => n2242, B2 => n694,
                           ZN => n4271);
   U2952 : AOI221_X1 port map( B1 => n697, B2 => n4598, C1 => n700, C2 => n4630
                           , A => n4272, ZN => n4265);
   U2953 : OAI22_X1 port map( A1 => n2244, A2 => n703, B1 => n2245, B2 => n706,
                           ZN => n4272);
   U2954 : NAND2_X1 port map( A1 => DATAIN(2), A2 => n264, ZN => n2217);
   U2955 : OAI21_X1 port map( B1 => n270, B2 => n4273, A => n710, ZN => n2987);
   U2956 : OAI221_X1 port map( B1 => n2247, B2 => n609, C1 => n276, C2 => n4274
                           , A => n4275, ZN => n2986);
   U2957 : OAI21_X1 port map( B1 => n4276, B2 => n4277, A => n610, ZN => n4275)
                           ;
   U2958 : NAND4_X1 port map( A1 => n4278, A2 => n4279, A3 => n4280, A4 => 
                           n4281, ZN => n4277);
   U2959 : AOI221_X1 port map( B1 => n613, B2 => n1060, C1 => n616, C2 => n1026
                           , A => n4282, ZN => n4281);
   U2960 : OAI22_X1 port map( A1 => n5045, A2 => n619, B1 => n5077, B2 => n622,
                           ZN => n4282);
   U2961 : AOI221_X1 port map( B1 => n625, B2 => n888, C1 => n628, C2 => n922, 
                           A => n4283, ZN => n4280);
   U2962 : OAI22_X1 port map( A1 => n5333, A2 => n631, B1 => n5301, B2 => n634,
                           ZN => n4283);
   U2963 : AOI221_X1 port map( B1 => n637, B2 => n2246, C1 => n640, C2 => n1309
                           , A => n4284, ZN => n4279);
   U2964 : OAI22_X1 port map( A1 => n4469, A2 => n643, B1 => n4501, B2 => n646,
                           ZN => n4284);
   U2965 : AOI221_X1 port map( B1 => n649, B2 => n1130, C1 => n652, C2 => n1096
                           , A => n4285, ZN => n4278);
   U2966 : OAI22_X1 port map( A1 => n4661, A2 => n655, B1 => n4693, B2 => n658,
                           ZN => n4285);
   U2967 : NAND4_X1 port map( A1 => n4286, A2 => n4287, A3 => n4288, A4 => 
                           n4289, ZN => n4276);
   U2968 : AOI221_X1 port map( B1 => n661, B2 => n4981, C1 => n664, C2 => n5013
                           , A => n4290, ZN => n4289);
   U2969 : OAI22_X1 port map( A1 => n2265, A2 => n667, B1 => n2266, B2 => n670,
                           ZN => n4290);
   U2970 : AOI221_X1 port map( B1 => n673, B2 => n5269, C1 => n676, C2 => n5237
                           , A => n4291, ZN => n4288);
   U2971 : OAI22_X1 port map( A1 => n2268, A2 => n679, B1 => n2269, B2 => n682,
                           ZN => n4291);
   U2972 : AOI221_X1 port map( B1 => n685, B2 => n4533, C1 => n688, C2 => n4565
                           , A => n4292, ZN => n4287);
   U2973 : OAI22_X1 port map( A1 => n2271, A2 => n691, B1 => n2272, B2 => n694,
                           ZN => n4292);
   U2974 : AOI221_X1 port map( B1 => n697, B2 => n4597, C1 => n700, C2 => n4629
                           , A => n4293, ZN => n4286);
   U2975 : OAI22_X1 port map( A1 => n2274, A2 => n703, B1 => n2275, B2 => n706,
                           ZN => n4293);
   U2976 : NAND2_X1 port map( A1 => DATAIN(1), A2 => n262, ZN => n2247);
   U2977 : OAI21_X1 port map( B1 => n270, B2 => n4294, A => n710, ZN => n2985);
   U2978 : OAI221_X1 port map( B1 => n2277, B2 => n609, C1 => n276, C2 => n4295
                           , A => n4296, ZN => n2984);
   U2979 : OAI21_X1 port map( B1 => n4297, B2 => n4298, A => n610, ZN => n4296)
                           ;
   U2980 : AND2_X1 port map( A1 => n609, A2 => n276, ZN => n2334);
   U2981 : NAND4_X1 port map( A1 => n4299, A2 => n4300, A3 => n4301, A4 => 
                           n4302, ZN => n4298);
   U2982 : AOI221_X1 port map( B1 => n613, B2 => n1061, C1 => n616, C2 => n1027
                           , A => n4303, ZN => n4302);
   U2983 : OAI22_X1 port map( A1 => n5044, A2 => n619, B1 => n5076, B2 => n622,
                           ZN => n4303);
   U2984 : NAND2_X1 port map( A1 => n4304, A2 => n4305, ZN => n2343);
   U2985 : NAND2_X1 port map( A1 => n4304, A2 => n4306, ZN => n2342);
   U2986 : AND2_X1 port map( A1 => n4307, A2 => n4305, ZN => n2340);
   U2987 : AND2_X1 port map( A1 => n4307, A2 => n4306, ZN => n2339);
   U2988 : AOI221_X1 port map( B1 => n625, B2 => n889, C1 => n628, C2 => n923, 
                           A => n4308, ZN => n4301);
   U2989 : OAI22_X1 port map( A1 => n5332, A2 => n631, B1 => n5300, B2 => n634,
                           ZN => n4308);
   U2990 : NAND2_X1 port map( A1 => n4304, A2 => n4309, ZN => n2348);
   U2991 : NAND2_X1 port map( A1 => n4304, A2 => n4310, ZN => n2347);
   U2992 : AND2_X1 port map( A1 => n4307, A2 => n4309, ZN => n2345);
   U2993 : AND2_X1 port map( A1 => n4307, A2 => n4310, ZN => n2344);
   U2994 : AOI221_X1 port map( B1 => n637, B2 => n2276, C1 => n640, C2 => n1310
                           , A => n4311, ZN => n4300);
   U2995 : OAI22_X1 port map( A1 => n4468, A2 => n643, B1 => n4500, B2 => n646,
                           ZN => n4311);
   U2996 : NAND2_X1 port map( A1 => n4312, A2 => n4313, ZN => n2353);
   U2997 : NAND2_X1 port map( A1 => n4314, A2 => n4313, ZN => n2352);
   U2998 : AND2_X1 port map( A1 => n4312, A2 => n4315, ZN => n2350);
   U2999 : AND2_X1 port map( A1 => n4314, A2 => n4315, ZN => n2349);
   U3000 : AOI221_X1 port map( B1 => n649, B2 => n1131, C1 => n652, C2 => n1097
                           , A => n4316, ZN => n4299);
   U3001 : OAI22_X1 port map( A1 => n4660, A2 => n655, B1 => n4692, B2 => n658,
                           ZN => n4316);
   U3002 : NAND2_X1 port map( A1 => n4317, A2 => n4307, ZN => n2358);
   U3003 : NAND2_X1 port map( A1 => n4318, A2 => n4307, ZN => n2357);
   U3004 : AND2_X1 port map( A1 => n4317, A2 => n4304, ZN => n2355);
   U3005 : AND2_X1 port map( A1 => n4318, A2 => n4304, ZN => n2354);
   U3006 : NAND4_X1 port map( A1 => n4319, A2 => n4320, A3 => n4321, A4 => 
                           n4322, ZN => n4297);
   U3007 : AOI221_X1 port map( B1 => n661, B2 => n4980, C1 => n664, C2 => n5012
                           , A => n4323, ZN => n4322);
   U3008 : OAI22_X1 port map( A1 => n2307, A2 => n667, B1 => n2308, B2 => n670,
                           ZN => n4323);
   U3009 : NAND2_X1 port map( A1 => n4315, A2 => n4305, ZN => n2367);
   U3010 : NAND2_X1 port map( A1 => n4315, A2 => n4306, ZN => n2366);
   U3011 : AND2_X1 port map( A1 => n4305, A2 => n4313, ZN => n2364);
   U3012 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(4), A3 => n4324, 
                           ZN => n4305);
   U3013 : AND2_X1 port map( A1 => n4313, A2 => n4306, ZN => n2363);
   U3014 : NOR3_X1 port map( A1 => n4325, A2 => ADD_RD1(4), A3 => n4324, ZN => 
                           n4306);
   U3015 : AOI221_X1 port map( B1 => n673, B2 => n5268, C1 => n676, C2 => n5236
                           , A => n4326, ZN => n4321);
   U3016 : OAI22_X1 port map( A1 => n2312, A2 => n679, B1 => n2313, B2 => n682,
                           ZN => n4326);
   U3017 : NAND2_X1 port map( A1 => n4309, A2 => n4315, ZN => n2372);
   U3018 : NAND2_X1 port map( A1 => n4310, A2 => n4315, ZN => n2371);
   U3019 : AND2_X1 port map( A1 => n4309, A2 => n4313, ZN => n2369);
   U3020 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => n4325, 
                           ZN => n4309);
   U3021 : AND2_X1 port map( A1 => n4310, A2 => n4313, ZN => n2368);
   U3022 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => 
                           ADD_RD1(0), ZN => n4310);
   U3023 : AOI221_X1 port map( B1 => n685, B2 => n4532, C1 => n688, C2 => n4564
                           , A => n4327, ZN => n4320);
   U3024 : OAI22_X1 port map( A1 => n2315, A2 => n691, B1 => n2316, B2 => n694,
                           ZN => n4327);
   U3025 : NAND2_X1 port map( A1 => n4307, A2 => n4312, ZN => n2377);
   U3026 : NAND2_X1 port map( A1 => n4307, A2 => n4314, ZN => n2376);
   U3027 : NOR2_X1 port map( A1 => n4328, A2 => ADD_RD1(1), ZN => n4307);
   U3028 : AND2_X1 port map( A1 => n4312, A2 => n4304, ZN => n2374);
   U3029 : NOR3_X1 port map( A1 => n4329, A2 => ADD_RD1(0), A3 => n4324, ZN => 
                           n4312);
   U3030 : AND2_X1 port map( A1 => n4304, A2 => n4314, ZN => n2373);
   U3031 : NOR3_X1 port map( A1 => n4329, A2 => n4325, A3 => n4324, ZN => n4314
                           );
   U3032 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n4304);
   U3033 : AOI221_X1 port map( B1 => n697, B2 => n4596, C1 => n700, C2 => n4628
                           , A => n4330, ZN => n4319);
   U3034 : OAI22_X1 port map( A1 => n2320, A2 => n703, B1 => n2321, B2 => n706,
                           ZN => n4330);
   U3035 : NAND2_X1 port map( A1 => n4317, A2 => n4313, ZN => n2382);
   U3036 : NAND2_X1 port map( A1 => n4318, A2 => n4313, ZN => n2381);
   U3037 : NOR2_X1 port map( A1 => n4331, A2 => ADD_RD1(2), ZN => n4313);
   U3038 : AND2_X1 port map( A1 => n4317, A2 => n4315, ZN => n2379);
   U3039 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(3), A3 => n4329, 
                           ZN => n4317);
   U3040 : AND2_X1 port map( A1 => n4318, A2 => n4315, ZN => n2378);
   U3041 : NOR2_X1 port map( A1 => n4328, A2 => n4331, ZN => n4315);
   U3042 : INV_X1 port map( A => ADD_RD1(1), ZN => n4331);
   U3043 : NOR3_X1 port map( A1 => n4325, A2 => ADD_RD1(3), A3 => n4329, ZN => 
                           n4318);
   U3044 : INV_X1 port map( A => ADD_RD1(0), ZN => n4325);
   U3045 : NAND4_X1 port map( A1 => n4332, A2 => n4333, A3 => n4334, A4 => 
                           n4335, ZN => n2329);
   U3046 : NOR4_X1 port map( A1 => n1064, A2 => n4336, A3 => n4337, A4 => n4338
                           , ZN => n4335);
   U3047 : XOR2_X1 port map( A => ADD_WR(1), B => ADD_RD1(1), Z => n4338);
   U3048 : XOR2_X1 port map( A => ADD_WR(0), B => ADD_RD1(0), Z => n4337);
   U3049 : INV_X1 port map( A => WR, ZN => n1064);
   U3050 : XOR2_X1 port map( A => n4324, B => ADD_WR(3), Z => n4334);
   U3051 : INV_X1 port map( A => ADD_RD1(3), ZN => n4324);
   U3052 : XOR2_X1 port map( A => ADD_WR(4), B => n4329, Z => n4333);
   U3053 : INV_X1 port map( A => ADD_RD1(4), ZN => n4329);
   U3054 : XOR2_X1 port map( A => n4328, B => ADD_WR(2), Z => n4332);
   U3055 : INV_X1 port map( A => ADD_RD1(2), ZN => n4328);
   U3056 : NAND2_X1 port map( A1 => DATAIN(0), A2 => n262, ZN => n2277);
   U3057 : OAI21_X1 port map( B1 => n267, B2 => n4339, A => n710, ZN => n2983);
   U3058 : OAI21_X1 port map( B1 => n747, B2 => n4336, A => n260, ZN => n2384);
   U3059 : INV_X1 port map( A => RD1, ZN => n4336);
   U3060 : INV_X1 port map( A => ENABLE, ZN => n747);
   U3061 : INV_X1 port map( A => RESET, ZN => n713);

end SYN_A;

library IEEE;

use IEEE.std_logic_1164.all;

use 
   work.CONV_PACK_windowedRegisterFile_size_word32_m_global5_n_in_out_local2_f_windows4_size_ext_addr4.all;

entity controUnit_f_windows6_size_windows3 is

   port( clock, reset, enable, call, ret, mmu_done : in std_logic;  fill, spill
         : out std_logic;  cwp_out : out std_logic_vector (2 downto 0));

end controUnit_f_windows6_size_windows3;

architecture SYN_behavioral of controUnit_f_windows6_size_windows3 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal cwp_out_2_port, cwp_out_1_port, cwp_out_0_port, currentState_2_port, 
      currentState_1_port, currentState_0_port, nextState_2_port, 
      nextState_1_port, nextState_0_port, canRestore_2_port, canRestore_1_port,
      canRestore_0_port, canSave_2_port, canSave_1_port, canSave_0_port, N106, 
      N108, N110, N112, N114, N116, N118, N120, N122, N124, N126, N130, N131, 
      N132, N144, N153, N154, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64 : std_logic;

begin
   cwp_out <= ( cwp_out_2_port, cwp_out_1_port, cwp_out_0_port );
   
   canSave_reg_0_inst : DLH_X1 port map( G => N153, D => N118, Q => 
                           canSave_0_port);
   canSave_reg_1_inst : DLH_X1 port map( G => N153, D => N120, Q => 
                           canSave_1_port);
   canSave_reg_2_inst : DLH_X1 port map( G => N153, D => N122, Q => 
                           canSave_2_port);
   nextState_reg_0_inst : DLH_X1 port map( G => enable, D => N130, Q => 
                           nextState_0_port);
   currentState_reg_0_inst : DFF_X1 port map( D => nextState_0_port, CK => 
                           clock, Q => currentState_0_port, QN => n14);
   nextState_reg_1_inst : DLH_X1 port map( G => enable, D => N131, Q => 
                           nextState_1_port);
   currentState_reg_1_inst : DFF_X1 port map( D => nextState_1_port, CK => 
                           clock, Q => currentState_1_port, QN => n30);
   canRestore_reg_1_inst : DLH_X1 port map( G => N153, D => N114, Q => 
                           canRestore_1_port);
   canRestore_reg_2_inst : DLH_X1 port map( G => N153, D => N116, Q => 
                           canRestore_2_port);
   nextState_reg_2_inst : DLH_X1 port map( G => enable, D => N132, Q => 
                           nextState_2_port);
   currentState_reg_2_inst : DFF_X1 port map( D => nextState_2_port, CK => 
                           clock, Q => currentState_2_port, QN => n6);
   fill_reg : DLH_X1 port map( G => N154, D => N124, Q => fill);
   canRestore_reg_0_inst : DLH_X1 port map( G => N153, D => N112, Q => 
                           canRestore_0_port);
   spill_reg : DLH_X1 port map( G => N144, D => N126, Q => spill);
   cwp_reg_0_inst : DLL_X1 port map( D => N106, GN => n16, Q => cwp_out_0_port)
                           ;
   cwp_reg_1_inst : DLL_X1 port map( D => N108, GN => n16, Q => cwp_out_1_port)
                           ;
   cwp_reg_2_inst : DLL_X1 port map( D => N110, GN => n16, Q => cwp_out_2_port)
                           ;
   U68 : XOR2_X1 port map( A => n36, B => canSave_2_port, Z => n34);
   U69 : XOR2_X1 port map( A => n45, B => canRestore_2_port, Z => n42);
   U70 : XOR2_X1 port map( A => canRestore_1_port, B => canRestore_0_port, Z =>
                           n47);
   U71 : NAND3_X1 port map( A1 => n27, A2 => n55, A3 => n53, ZN => n54);
   U72 : NAND3_X1 port map( A1 => n24, A2 => n59, A3 => call, ZN => n52);
   U73 : NAND3_X1 port map( A1 => n51, A2 => n60, A3 => cwp_out_0_port, ZN => 
                           n59);
   U74 : XOR2_X1 port map( A => cwp_out_2_port, B => n63, Z => n49);
   U75 : XOR2_X1 port map( A => cwp_out_1_port, B => cwp_out_0_port, Z => n60);
   U3 : NOR3_X1 port map( A1 => currentState_0_port, A2 => currentState_2_port,
                           A3 => n30, ZN => N126);
   U4 : NOR3_X1 port map( A1 => n24, A2 => N124, A3 => N126, ZN => n41);
   U5 : NOR2_X1 port map( A1 => N126, A2 => n27, ZN => n33);
   U6 : AOI22_X1 port map( A1 => n20, A2 => N126, B1 => n9, B2 => N124, ZN => 
                           n15);
   U7 : OAI21_X1 port map( B1 => n15, B2 => n8, A => n16, ZN => N153);
   U8 : INV_X1 port map( A => n10, ZN => n35);
   U9 : INV_X1 port map( A => n56, ZN => n27);
   U10 : OAI21_X1 port map( B1 => n52, B2 => n53, A => n54, ZN => N108);
   U11 : INV_X1 port map( A => n52, ZN => n50);
   U12 : NAND2_X1 port map( A1 => n53, A2 => n49, ZN => n58);
   U13 : INV_X1 port map( A => n60, ZN => n53);
   U14 : INV_X1 port map( A => n38, ZN => n37);
   U15 : INV_X1 port map( A => n48, ZN => N110);
   U16 : AOI221_X1 port map( B1 => n49, B2 => n27, C1 => n50, C2 => n51, A => 
                           n10, ZN => n48);
   U17 : NOR3_X1 port map( A1 => currentState_1_port, A2 => currentState_2_port
                           , A3 => currentState_0_port, ZN => n10);
   U18 : NOR3_X1 port map( A1 => n14, A2 => currentState_2_port, A3 => n30, ZN 
                           => N124);
   U19 : NOR3_X1 port map( A1 => currentState_1_port, A2 => currentState_2_port
                           , A3 => n14, ZN => n24);
   U20 : NOR2_X1 port map( A1 => cwp_out_0_port, A2 => cwp_out_1_port, ZN => 
                           n63);
   U21 : AOI21_X1 port map( B1 => n24, B2 => call, A => N124, ZN => n31);
   U22 : NOR2_X1 port map( A1 => n37, A2 => canSave_2_port, ZN => n20);
   U23 : AOI22_X1 port map( A1 => enable, A2 => N131, B1 => n17, B2 => n10, ZN 
                           => n16);
   U24 : INV_X1 port map( A => n8, ZN => n17);
   U25 : NOR2_X1 port map( A1 => n44, A2 => canRestore_2_port, ZN => n9);
   U26 : OAI221_X1 port map( B1 => n31, B2 => n32, C1 => n33, C2 => n34, A => 
                           n35, ZN => N122);
   U27 : AOI21_X1 port map( B1 => canSave_2_port, B2 => n37, A => n20, ZN => 
                           n32);
   U28 : NAND2_X1 port map( A1 => canSave_1_port, A2 => canSave_0_port, ZN => 
                           n36);
   U29 : OAI221_X1 port map( B1 => n33, B2 => n39, C1 => n31, C2 => n40, A => 
                           n35, ZN => N120);
   U30 : INV_X1 port map( A => n40, ZN => n39);
   U31 : AOI21_X1 port map( B1 => canSave_0_port, B2 => canSave_1_port, A => 
                           n38, ZN => n40);
   U32 : OAI221_X1 port map( B1 => n56, B2 => n55, C1 => cwp_out_0_port, C2 => 
                           n57, A => n35, ZN => N106);
   U33 : AOI21_X1 port map( B1 => n27, B2 => n58, A => n50, ZN => n57);
   U34 : OAI22_X1 port map( A1 => n31, A2 => n42, B1 => n33, B2 => n43, ZN => 
                           N116);
   U35 : AOI21_X1 port map( B1 => canRestore_2_port, B2 => n44, A => n9, ZN => 
                           n43);
   U36 : NAND2_X1 port map( A1 => canRestore_1_port, A2 => canRestore_0_port, 
                           ZN => n45);
   U37 : OAI22_X1 port map( A1 => n31, A2 => n46, B1 => n33, B2 => n47, ZN => 
                           N114);
   U38 : INV_X1 port map( A => n47, ZN => n46);
   U39 : NOR2_X1 port map( A1 => canSave_1_port, A2 => canSave_0_port, ZN => 
                           n38);
   U40 : XNOR2_X1 port map( A => n61, B => cwp_out_2_port, ZN => n51);
   U41 : NAND2_X1 port map( A1 => cwp_out_0_port, A2 => cwp_out_1_port, ZN => 
                           n61);
   U42 : NAND2_X1 port map( A1 => n24, A2 => n64, ZN => n56);
   U43 : INV_X1 port map( A => call, ZN => n64);
   U44 : NAND2_X1 port map( A1 => currentState_2_port, A2 => n30, ZN => n13);
   U45 : AOI21_X1 port map( B1 => n12, B2 => n14, A => n13, ZN => n29);
   U46 : NAND2_X1 port map( A1 => enable, A2 => n19, ZN => n8);
   U47 : AOI21_X1 port map( B1 => n25, B2 => n26, A => reset, ZN => N130);
   U48 : AOI21_X1 port map( B1 => N126, B2 => n28, A => n29, ZN => n25);
   U49 : NOR3_X1 port map( A1 => N124, A2 => n10, A3 => n27, ZN => n26);
   U50 : INV_X1 port map( A => n20, ZN => n28);
   U51 : INV_X1 port map( A => mmu_done, ZN => n12);
   U52 : NAND2_X1 port map( A1 => n62, A2 => cwp_out_0_port, ZN => n55);
   U53 : INV_X1 port map( A => n58, ZN => n62);
   U54 : NOR2_X1 port map( A1 => n18, A2 => n8, ZN => N144);
   U55 : AOI211_X1 port map( C1 => N126, C2 => n20, A => n10, B => n21, ZN => 
                           n18);
   U56 : NOR3_X1 port map( A1 => n12, A2 => currentState_0_port, A3 => n13, ZN 
                           => n21);
   U57 : NOR2_X1 port map( A1 => n7, A2 => n8, ZN => N154);
   U58 : AOI211_X1 port map( C1 => N124, C2 => n9, A => n10, B => n11, ZN => n7
                           );
   U59 : NOR3_X1 port map( A1 => n12, A2 => n13, A3 => n14, ZN => n11);
   U60 : INV_X1 port map( A => reset, ZN => n19);
   U61 : NOR2_X1 port map( A1 => canSave_0_port, A2 => n41, ZN => N118);
   U62 : NOR2_X1 port map( A1 => canRestore_0_port, A2 => n41, ZN => N112);
   U63 : OR2_X1 port map( A1 => canRestore_1_port, A2 => canRestore_0_port, ZN 
                           => n44);
   U64 : INV_X1 port map( A => n23, ZN => N131);
   U65 : OAI211_X1 port map( C1 => call, C2 => ret, A => n19, B => n24, ZN => 
                           n23);
   U66 : AND2_X1 port map( A1 => n19, A2 => n22, ZN => N132);
   U67 : OAI21_X1 port map( B1 => n13, B2 => mmu_done, A => n15, ZN => n22);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use 
   work.CONV_PACK_windowedRegisterFile_size_word32_m_global5_n_in_out_local2_f_windows4_size_ext_addr4.all;

entity 
   windowedRegisterFile_size_word32_m_global5_n_in_out_local2_f_windows4_size_ext_addr4 
   is

   port( data_in_write : in std_logic_vector (31 downto 0);  addr_write, 
         addr_read_one, addr_read_two : in std_logic_vector (3 downto 0);  
         data_out_port_one, data_out_port_two : out std_logic_vector (31 downto
         0);  fill, spill : out std_logic;  call, ret, mmu_done, clock, reset, 
         enable, read_en_one, read_en_two, write_en : in std_logic);

end 
   windowedRegisterFile_size_word32_m_global5_n_in_out_local2_f_windows4_size_ext_addr4;

architecture SYN_structural of 
   windowedRegisterFile_size_word32_m_global5_n_in_out_local2_f_windows4_size_ext_addr4 
   is

   component register_file_nBitsData32_nBitsAddr5
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component controUnit_f_windows6_size_windows3
      port( clock, reset, enable, call, ret, mmu_done : in std_logic;  fill, 
            spill : out std_logic;  cwp_out : out std_logic_vector (2 downto 0)
            );
   end component;
   
   component addressesGenerator
      port( addr_read_one_in, addr_read_two_in, addr_write_in : in 
            std_logic_vector (3 downto 0);  cwp_in : in std_logic_vector (2 
            downto 0);  addr_read_one_out, addr_read_two_out, addr_write_out : 
            out std_logic_vector (4 downto 0));
   end component;
   
   signal cwp_s_1_port, cwp_s_0_port, addr_read_one_s_4_port, 
      addr_read_one_s_3_port, addr_read_one_s_2_port, addr_read_one_s_1_port, 
      addr_read_one_s_0_port, addr_read_two_s_4_port, addr_read_two_s_3_port, 
      addr_read_two_s_2_port, addr_read_two_s_1_port, addr_read_two_s_0_port, 
      addr_write_s_4_port, addr_write_s_3_port, addr_write_s_2_port, 
      addr_write_s_1_port, addr_write_s_0_port, n1, n_1000 : std_logic;

begin
   
   m_AD : addressesGenerator port map( addr_read_one_in(3) => addr_read_one(3),
                           addr_read_one_in(2) => addr_read_one(2), 
                           addr_read_one_in(1) => addr_read_one(1), 
                           addr_read_one_in(0) => addr_read_one(0), 
                           addr_read_two_in(3) => addr_read_two(3), 
                           addr_read_two_in(2) => addr_read_two(2), 
                           addr_read_two_in(1) => addr_read_two(1), 
                           addr_read_two_in(0) => addr_read_two(0), 
                           addr_write_in(3) => addr_write(3), addr_write_in(2) 
                           => addr_write(2), addr_write_in(1) => addr_write(1),
                           addr_write_in(0) => addr_write(0), cwp_in(2) => n1, 
                           cwp_in(1) => cwp_s_1_port, cwp_in(0) => cwp_s_0_port
                           , addr_read_one_out(4) => addr_read_one_s_4_port, 
                           addr_read_one_out(3) => addr_read_one_s_3_port, 
                           addr_read_one_out(2) => addr_read_one_s_2_port, 
                           addr_read_one_out(1) => addr_read_one_s_1_port, 
                           addr_read_one_out(0) => addr_read_one_s_0_port, 
                           addr_read_two_out(4) => addr_read_two_s_4_port, 
                           addr_read_two_out(3) => addr_read_two_s_3_port, 
                           addr_read_two_out(2) => addr_read_two_s_2_port, 
                           addr_read_two_out(1) => addr_read_two_s_1_port, 
                           addr_read_two_out(0) => addr_read_two_s_0_port, 
                           addr_write_out(4) => addr_write_s_4_port, 
                           addr_write_out(3) => addr_write_s_3_port, 
                           addr_write_out(2) => addr_write_s_2_port, 
                           addr_write_out(1) => addr_write_s_1_port, 
                           addr_write_out(0) => addr_write_s_0_port);
   m_CU : controUnit_f_windows6_size_windows3 port map( clock => clock, reset 
                           => reset, enable => enable, call => call, ret => ret
                           , mmu_done => mmu_done, fill => fill, spill => spill
                           , cwp_out(2) => n_1000, cwp_out(1) => cwp_s_1_port, 
                           cwp_out(0) => cwp_s_0_port);
   m_RF : register_file_nBitsData32_nBitsAddr5 port map( CLK => clock, RESET =>
                           reset, ENABLE => enable, RD1 => read_en_one, RD2 => 
                           read_en_two, WR => write_en, ADD_WR(4) => 
                           addr_write_s_4_port, ADD_WR(3) => 
                           addr_write_s_3_port, ADD_WR(2) => 
                           addr_write_s_2_port, ADD_WR(1) => 
                           addr_write_s_1_port, ADD_WR(0) => 
                           addr_write_s_0_port, ADD_RD1(4) => 
                           addr_read_one_s_4_port, ADD_RD1(3) => 
                           addr_read_one_s_3_port, ADD_RD1(2) => 
                           addr_read_one_s_2_port, ADD_RD1(1) => 
                           addr_read_one_s_1_port, ADD_RD1(0) => 
                           addr_read_one_s_0_port, ADD_RD2(4) => 
                           addr_read_two_s_4_port, ADD_RD2(3) => 
                           addr_read_two_s_3_port, ADD_RD2(2) => 
                           addr_read_two_s_2_port, ADD_RD2(1) => 
                           addr_read_two_s_1_port, ADD_RD2(0) => 
                           addr_read_two_s_0_port, DATAIN(31) => 
                           data_in_write(31), DATAIN(30) => data_in_write(30), 
                           DATAIN(29) => data_in_write(29), DATAIN(28) => 
                           data_in_write(28), DATAIN(27) => data_in_write(27), 
                           DATAIN(26) => data_in_write(26), DATAIN(25) => 
                           data_in_write(25), DATAIN(24) => data_in_write(24), 
                           DATAIN(23) => data_in_write(23), DATAIN(22) => 
                           data_in_write(22), DATAIN(21) => data_in_write(21), 
                           DATAIN(20) => data_in_write(20), DATAIN(19) => 
                           data_in_write(19), DATAIN(18) => data_in_write(18), 
                           DATAIN(17) => data_in_write(17), DATAIN(16) => 
                           data_in_write(16), DATAIN(15) => data_in_write(15), 
                           DATAIN(14) => data_in_write(14), DATAIN(13) => 
                           data_in_write(13), DATAIN(12) => data_in_write(12), 
                           DATAIN(11) => data_in_write(11), DATAIN(10) => 
                           data_in_write(10), DATAIN(9) => data_in_write(9), 
                           DATAIN(8) => data_in_write(8), DATAIN(7) => 
                           data_in_write(7), DATAIN(6) => data_in_write(6), 
                           DATAIN(5) => data_in_write(5), DATAIN(4) => 
                           data_in_write(4), DATAIN(3) => data_in_write(3), 
                           DATAIN(2) => data_in_write(2), DATAIN(1) => 
                           data_in_write(1), DATAIN(0) => data_in_write(0), 
                           OUT1(31) => data_out_port_one(31), OUT1(30) => 
                           data_out_port_one(30), OUT1(29) => 
                           data_out_port_one(29), OUT1(28) => 
                           data_out_port_one(28), OUT1(27) => 
                           data_out_port_one(27), OUT1(26) => 
                           data_out_port_one(26), OUT1(25) => 
                           data_out_port_one(25), OUT1(24) => 
                           data_out_port_one(24), OUT1(23) => 
                           data_out_port_one(23), OUT1(22) => 
                           data_out_port_one(22), OUT1(21) => 
                           data_out_port_one(21), OUT1(20) => 
                           data_out_port_one(20), OUT1(19) => 
                           data_out_port_one(19), OUT1(18) => 
                           data_out_port_one(18), OUT1(17) => 
                           data_out_port_one(17), OUT1(16) => 
                           data_out_port_one(16), OUT1(15) => 
                           data_out_port_one(15), OUT1(14) => 
                           data_out_port_one(14), OUT1(13) => 
                           data_out_port_one(13), OUT1(12) => 
                           data_out_port_one(12), OUT1(11) => 
                           data_out_port_one(11), OUT1(10) => 
                           data_out_port_one(10), OUT1(9) => 
                           data_out_port_one(9), OUT1(8) => 
                           data_out_port_one(8), OUT1(7) => 
                           data_out_port_one(7), OUT1(6) => 
                           data_out_port_one(6), OUT1(5) => 
                           data_out_port_one(5), OUT1(4) => 
                           data_out_port_one(4), OUT1(3) => 
                           data_out_port_one(3), OUT1(2) => 
                           data_out_port_one(2), OUT1(1) => 
                           data_out_port_one(1), OUT1(0) => 
                           data_out_port_one(0), OUT2(31) => 
                           data_out_port_two(31), OUT2(30) => 
                           data_out_port_two(30), OUT2(29) => 
                           data_out_port_two(29), OUT2(28) => 
                           data_out_port_two(28), OUT2(27) => 
                           data_out_port_two(27), OUT2(26) => 
                           data_out_port_two(26), OUT2(25) => 
                           data_out_port_two(25), OUT2(24) => 
                           data_out_port_two(24), OUT2(23) => 
                           data_out_port_two(23), OUT2(22) => 
                           data_out_port_two(22), OUT2(21) => 
                           data_out_port_two(21), OUT2(20) => 
                           data_out_port_two(20), OUT2(19) => 
                           data_out_port_two(19), OUT2(18) => 
                           data_out_port_two(18), OUT2(17) => 
                           data_out_port_two(17), OUT2(16) => 
                           data_out_port_two(16), OUT2(15) => 
                           data_out_port_two(15), OUT2(14) => 
                           data_out_port_two(14), OUT2(13) => 
                           data_out_port_two(13), OUT2(12) => 
                           data_out_port_two(12), OUT2(11) => 
                           data_out_port_two(11), OUT2(10) => 
                           data_out_port_two(10), OUT2(9) => 
                           data_out_port_two(9), OUT2(8) => 
                           data_out_port_two(8), OUT2(7) => 
                           data_out_port_two(7), OUT2(6) => 
                           data_out_port_two(6), OUT2(5) => 
                           data_out_port_two(5), OUT2(4) => 
                           data_out_port_two(4), OUT2(3) => 
                           data_out_port_two(3), OUT2(2) => 
                           data_out_port_two(2), OUT2(1) => 
                           data_out_port_two(1), OUT2(0) => 
                           data_out_port_two(0));
   n1 <= '0';

end SYN_structural;
