
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_register_file_nBitsData64_nBitsAddr5 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_register_file_nBitsData64_nBitsAddr5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_register_file_nBitsData64_nBitsAddr5.all;

entity register_file_nBitsData64_nBitsAddr5 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector (63
         downto 0));

end register_file_nBitsData64_nBitsAddr5;

architecture SYN_A of register_file_nBitsData64_nBitsAddr5 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component TINV_X1
      port( I, EN : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5130, n5132, n5134, n5136, n5138, n5140, n5142, n5144, n5146, n5148,
      n5150, n5152, n5154, n5156, n5158, n5160, n5162, n5164, n5166, n5168, 
      n5170, n5172, n5174, n5176, n5178, n5180, n5182, n5184, n5186, n5188, 
      n5190, n5192, n5194, n5196, n5198, n5200, n5202, n5204, n5206, n5208, 
      n5210, n5212, n5214, n5216, n5218, n5220, n5222, n5224, n5226, n5228, 
      n5230, n5232, n5234, n5236, n5238, n5240, n5242, n5244, n5246, n5248, 
      n5250, n5252, n5254, n5256, n5258, n5260, n5262, n5264, n5266, n5268, 
      n5270, n5272, n5274, n5276, n5278, n5280, n5282, n5284, n5286, n5288, 
      n5290, n5292, n5294, n5296, n5298, n5300, n5302, n5304, n5306, n5308, 
      n5310, n5312, n5314, n5316, n5318, n5320, n5322, n5324, n5326, n5328, 
      n5330, n5332, n5334, n5336, n5338, n5340, n5342, n5344, n5346, n5348, 
      n5350, n5352, n5354, n5356, n5358, n5360, n5362, n5364, n5366, n5368, 
      n5370, n5372, n5374, n5376, n5378, n5380, n5382, n5384, n5641, n5642, 
      n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, 
      n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, 
      n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, 
      n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, 
      n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, 
      n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, 
      n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, 
      n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, 
      n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, 
      n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, 
      n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, 
      n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, 
      n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, 
      n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, 
      n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, 
      n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, 
      n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, 
      n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, 
      n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, 
      n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, 
      n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, 
      n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, 
      n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, 
      n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, 
      n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, 
      n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, 
      n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, 
      n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, 
      n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, 
      n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, 
      n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, 
      n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, 
      n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, 
      n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, 
      n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, 
      n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, 
      n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, 
      n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, 
      n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, 
      n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, 
      n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, 
      n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, 
      n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, 
      n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, 
      n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, 
      n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, 
      n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, 
      n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, 
      n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, 
      n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, 
      n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, 
      n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, 
      n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, 
      n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, 
      n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, 
      n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, 
      n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, 
      n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, 
      n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, 
      n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, 
      n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, 
      n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, 
      n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, 
      n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, 
      n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, 
      n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, 
      n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, 
      n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, 
      n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, 
      n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, 
      n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, 
      n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, 
      n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, 
      n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, 
      n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, 
      n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, 
      n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, 
      n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, 
      n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, 
      n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, 
      n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, 
      n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, 
      n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, 
      n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, 
      n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, 
      n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, 
      n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, 
      n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, 
      n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, 
      n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, 
      n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, 
      n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, 
      n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, 
      n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, 
      n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, 
      n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, 
      n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, 
      n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, 
      n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, 
      n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, 
      n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, 
      n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, 
      n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, 
      n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, 
      n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, 
      n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, 
      n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, 
      n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, 
      n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, 
      n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, 
      n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, 
      n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, 
      n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, 
      n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, 
      n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, 
      n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, 
      n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, 
      n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, 
      n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, 
      n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, 
      n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, 
      n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, 
      n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, 
      n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, 
      n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, 
      n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, 
      n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, 
      n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, 
      n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, 
      n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, 
      n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, 
      n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, 
      n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, 
      n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, 
      n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, 
      n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, 
      n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, 
      n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, 
      n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, 
      n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, 
      n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, 
      n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, 
      n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, 
      n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, 
      n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, 
      n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, 
      n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, 
      n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, 
      n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, 
      n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, 
      n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, 
      n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, 
      n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, 
      n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, 
      n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, 
      n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, 
      n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, 
      n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, 
      n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, 
      n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, 
      n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, 
      n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, 
      n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, 
      n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, 
      n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, 
      n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, 
      n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, 
      n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, 
      n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, 
      n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, 
      n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, 
      n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, 
      n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, 
      n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, 
      n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, 
      n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, 
      n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, 
      n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, 
      n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, 
      n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, 
      n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, 
      n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, 
      n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, 
      n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, 
      n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, 
      n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, 
      n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, 
      n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, 
      n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, 
      n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, 
      n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, 
      n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, 
      n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, 
      n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, 
      n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, 
      n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, 
      n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, 
      n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, 
      n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, 
      n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, 
      n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, 
      n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, 
      n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, 
      n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, 
      n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, 
      n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, 
      n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, 
      n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, 
      n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, 
      n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, 
      n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, 
      n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, 
      n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, 
      n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, 
      n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, 
      n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, 
      n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, 
      n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, 
      n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, 
      n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, 
      n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, 
      n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, 
      n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, 
      n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, 
      n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, 
      n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, 
      n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, 
      n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, 
      n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, 
      n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, 
      n7943, n7944, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, 
      n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, 
      n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, 
      n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, 
      n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, 
      n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, 
      n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, 
      n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, 
      n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, 
      n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, 
      n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, 
      n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, 
      n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, 
      n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, 
      n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, 
      n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, 
      n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, 
      n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, 
      n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, 
      n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, 
      n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, 
      n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, 
      n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, 
      n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, 
      n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, 
      n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, 
      n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, 
      n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, 
      n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, 
      n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, 
      n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, 
      n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, 
      n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, 
      n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, 
      n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, 
      n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, 
      n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, 
      n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, 
      n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, 
      n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, 
      n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, 
      n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, 
      n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, 
      n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, 
      n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, 
      n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, 
      n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, 
      n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, 
      n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, 
      n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, 
      n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, 
      n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, 
      n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, 
      n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, 
      n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, 
      n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, 
      n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, 
      n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, 
      n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, 
      n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, 
      n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, 
      n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, 
      n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, 
      n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, 
      n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, 
      n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, 
      n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, 
      n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, 
      n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, 
      n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, 
      n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, 
      n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, 
      n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, 
      n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, 
      n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, 
      n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, 
      n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, 
      n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, 
      n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, 
      n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, 
      n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, 
      n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, 
      n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, 
      n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, 
      n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, 
      n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, 
      n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, 
      n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, 
      n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, 
      n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, 
      n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, 
      n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, 
      n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, 
      n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, 
      n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, 
      n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, 
      n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, 
      n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, 
      n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, 
      n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, 
      n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, 
      n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, 
      n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, 
      n9997, n9998, n9999, n10761, n10762, n10763, n10764, n10765, n10766, 
      n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, 
      n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, 
      n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, 
      n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, 
      n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, 
      n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, 
      n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, 
      n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, 
      n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, 
      n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, 
      n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, 
      n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, 
      n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, 
      n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, 
      n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, 
      n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, 
      n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, 
      n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, 
      n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, 
      n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, 
      n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, 
      n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, 
      n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, 
      n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, 
      n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, 
      n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, 
      n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, 
      n11010, n11011, n11012, n11013, n11014, n11015, n11016, n13909, n13910, 
      n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919, 
      n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928, 
      n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937, 
      n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946, 
      n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955, 
      n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964, 
      n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13985, 
      n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994, 
      n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, 
      n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012, 
      n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021, 
      n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030, 
      n14031, n14032, n14033, n14034, n14035, n14036, n14549, n14550, n14551, 
      n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, 
      n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, 
      n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578, 
      n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, 
      n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596, 
      n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605, 
      n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14625, n14626, 
      n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635, 
      n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644, 
      n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653, 
      n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662, 
      n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671, 
      n14672, n14673, n14674, n14675, n14676, n15061, n15062, n15063, n15064, 
      n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073, 
      n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082, 
      n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091, 
      n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100, 
      n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109, 
      n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118, 
      n15119, n15120, n15121, n15122, n15123, n15124, n15136, n15137, n15138, 
      n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147, 
      n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156, 
      n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165, 
      n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174, 
      n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183, 
      n15184, n15185, n15186, n15187, n15188, n15445, n15446, n15447, n15448, 
      n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457, 
      n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466, 
      n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475, 
      n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484, 
      n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493, 
      n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502, 
      n15503, n15504, n15505, n15506, n15507, n15508, n15520, n15521, n15522, 
      n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531, 
      n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540, 
      n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549, 
      n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558, 
      n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567, 
      n15568, n15569, n15570, n15571, n15572, n15701, n15702, n15703, n15704, 
      n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713, 
      n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722, 
      n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731, 
      n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740, 
      n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749, 
      n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758, 
      n15759, n15760, n15761, n15762, n15763, n15764, n15776, n15777, n15778, 
      n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787, 
      n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796, 
      n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805, 
      n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814, 
      n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823, 
      n15824, n15825, n15826, n15827, n15828, n17772, n17774, n17775, n17776, 
      n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785, 
      n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794, 
      n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803, 
      n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812, 
      n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821, 
      n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830, 
      n17831, n17832, n17833, n17834, n17835, n17836, n18059, n18061, n18062, 
      n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071, 
      n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080, 
      n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089, 
      n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098, 
      n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107, 
      n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116, 
      n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18126, n18128, 
      n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137, 
      n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146, 
      n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155, 
      n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164, 
      n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173, 
      n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182, 
      n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18192, 
      n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202, 
      n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211, 
      n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220, 
      n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229, 
      n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238, 
      n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247, 
      n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256, 
      n18259, n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268, 
      n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277, 
      n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286, 
      n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295, 
      n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304, 
      n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313, 
      n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322, 
      n18323, n21795, n21796, n21797, n21798, n21799, n21800, n21801, n21802, 
      n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811, 
      n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820, 
      n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828, n21829, 
      n21830, n21831, n21832, n21833, n21834, n21835, n21836, n21837, n21838, 
      n21839, n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847, 
      n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856, 
      n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865, 
      n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21874, 
      n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883, 
      n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892, 
      n21893, n21894, n21895, n21896, n21897, n21898, n21899, n21900, n21901, 
      n21902, n21903, n21904, n21905, n21906, n21907, n21908, n21909, n21910, 
      n21911, n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919, 
      n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928, 
      n21929, n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937, 
      n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945, n21946, 
      n21947, n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955, 
      n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964, 
      n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972, n21973, 
      n21974, n21975, n21976, n21977, n21978, n21979, n21980, n21981, n21982, 
      n21983, n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991, 
      n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999, n22000, 
      n22001, n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009, 
      n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017, n22018, 
      n22019, n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027, 
      n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036, 
      n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044, n22045, 
      n22046, n22047, n22048, n22049, n22050, n22051, n22052, n22053, n22054, 
      n22055, n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063, 
      n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071, n22072, 
      n22073, n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081, 
      n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090, 
      n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099, 
      n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107, n22108, 
      n22109, n22110, n22111, n22112, n22113, n22114, n22179, n22180, n22181, 
      n22182, n22183, n22184, n22185, n22186, n22187, n22188, n22189, n22190, 
      n22191, n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199, 
      n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207, n22208, 
      n22209, n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217, 
      n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225, n22226, 
      n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235, 
      n22236, n22237, n22238, n22239, n22240, n22241, n22242, n25150, n25151, 
      n25152, n25153, n25154, n25155, n25156, n25157, n25158, n25159, n25160, 
      n25161, n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169, 
      n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177, n25178, 
      n25179, n25180, n25181, n25182, n25183, n25184, n25185, n25186, n25187, 
      n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195, n25196, 
      n25197, n25198, n25199, n25200, n25201, n25202, n25203, n25204, n25205, 
      n25206, n25207, n25208, n25209, n25210, n25211, n25212, n25213, n25214, 
      n25215, n25216, n25217, n25218, n25219, n25220, n25221, n25222, n25223, 
      n25224, n25225, n25226, n25227, n25228, n25229, n25230, n25231, n25232, 
      n25233, n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241, 
      n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249, n25250, 
      n25251, n25252, n25253, n25254, n25255, n25256, n25257, n25258, n25259, 
      n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267, n25268, 
      n25269, n25270, n25271, n25272, n25273, n25274, n25275, n25276, n25277, 
      n25278, n25279, n25280, n25281, n25282, n25283, n25284, n25285, n25286, 
      n25287, n25288, n25289, n25290, n25291, n25292, n25293, n25294, n25295, 
      n25296, n25297, n25298, n25299, n25300, n25301, n25302, n25303, n25304, 
      n25305, n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313, 
      n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321, n25322, 
      n25323, n25324, n25325, n25326, n25327, n25328, n25329, n25330, n25331, 
      n25332, n25333, n25334, n25335, n25336, n25337, n25338, n25339, n25340, 
      n25341, n25342, n25343, n25344, n25345, n25346, n25347, n25348, n25349, 
      n25350, n25351, n25352, n25353, n25354, n25355, n25356, n25357, n25358, 
      n25359, n25360, n25361, n25362, n25363, n25364, n25365, n25366, n25367, 
      n25368, n25369, n25370, n25371, n25372, n25373, n25374, n25375, n25376, 
      n25377, n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385, 
      n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393, n25394, 
      n25395, n25396, n25397, n25398, n25399, n25400, n25401, n25402, n25403, 
      n25404, n25405, n25406, n25407, n25408, n25409, n25410, n25411, n25412, 
      n25413, n25414, n25415, n25416, n25417, n25418, n25419, n25420, n25421, 
      n25422, n25423, n25424, n25425, n25426, n25427, n25428, n25429, n25430, 
      n25431, n25432, n25433, n25434, n25435, n25436, n25437, n25438, n25439, 
      n25440, n25441, n25442, n25443, n25444, n25445, n25446, n25447, n25448, 
      n25449, n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457, 
      n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465, n25466, 
      n25467, n25468, n25469, n25470, n25471, n25472, n25473, n25474, n25475, 
      n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483, n25484, 
      n25485, n25486, n25487, n25488, n25489, n25490, n25491, n25492, n25493, 
      n25494, n25495, n25496, n25497, n25498, n25499, n25500, n25501, n25502, 
      n25503, n25504, n25505, n25506, n25507, n25508, n25509, n25510, n25511, 
      n25512, n25513, n25514, n25515, n25516, n25517, n25518, n25519, n25520, 
      n25521, n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529, 
      n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537, n25538, 
      n25539, n25540, n25541, n25542, n25543, n25544, n25545, n25546, n25547, 
      n25548, n25549, n25550, n25551, n25552, n25553, n25554, n25555, n25556, 
      n25557, n25558, n25559, n25560, n25561, n25562, n25563, n25564, n25565, 
      n25566, n25567, n25568, n25569, n25570, n25571, n25572, n25573, n25574, 
      n25575, n25576, n25577, n25578, n25579, n25580, n25581, n25582, n25583, 
      n25584, n25585, n25586, n25587, n25588, n25589, n25590, n25591, n25592, 
      n25593, n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601, 
      n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609, n25610, 
      n25611, n25612, n25613, n25614, n25615, n25616, n25617, n25618, n25619, 
      n25620, n25621, n25622, n25623, n25624, n25625, n25626, n25627, n25628, 
      n25629, n25630, n25631, n25632, n25633, n25634, n25635, n25636, n25637, 
      n25638, n25639, n25640, n25641, n25642, n25643, n25644, n25645, n25646, 
      n25647, n25648, n25649, n25650, n25651, n25652, n25653, n25654, n25655, 
      n25656, n25657, n25658, n25659, n25660, n25661, n25662, n25663, n25664, 
      n25665, n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673, 
      n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681, n25682, 
      n25683, n25684, n25685, n25686, n25687, n25688, n25689, n25690, n25691, 
      n25692, n25693, n25694, n25695, n25696, n25697, n25698, n25699, n25700, 
      n25701, n25702, n25703, n25704, n25705, n25706, n25707, n25708, n25709, 
      n25710, n25711, n25712, n25713, n25714, n25715, n25716, n25717, n25718, 
      n25719, n25720, n25721, n25722, n25723, n25724, n25725, n25726, n25727, 
      n25728, n25729, n25730, n25731, n25732, n25733, n25734, n25735, n25736, 
      n25737, n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745, 
      n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753, n25754, 
      n25755, n25756, n25757, n25758, n25759, n25760, n25761, n25762, n25763, 
      n25764, n25765, n25766, n25767, n25768, n25769, n25770, n25771, n25772, 
      n25773, n25774, n25775, n25776, n25777, n25778, n25779, n25780, n25781, 
      n25782, n25783, n25784, n25785, n25786, n25787, n25788, n25789, n25790, 
      n25791, n25792, n25793, n25794, n25795, n25796, n25797, n25798, n25799, 
      n25800, n25801, n25802, n25803, n25804, n25805, n25806, n25807, n25808, 
      n25809, n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817, 
      n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825, n25826, 
      n25827, n25828, n25829, n25830, n25831, n25832, n25833, n25834, n25835, 
      n25836, n25837, n25838, n25839, n25840, n25841, n25842, n25843, n25844, 
      n25845, n25846, n25847, n25848, n25849, n25850, n25851, n25852, n25853, 
      n25854, n25855, n25856, n25857, n25858, n25859, n25860, n25861, n25862, 
      n25863, n25864, n25865, n25866, n25867, n25868, n25869, n25870, n25871, 
      n25872, n25873, n25874, n25875, n25876, n25877, n25878, n25879, n25880, 
      n25881, n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889, 
      n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897, n25898, 
      n25899, n25900, n25901, n25902, n25903, n25904, n25905, n25906, n25907, 
      n25908, n25909, n25910, n25911, n25912, n25913, n25914, n25915, n25916, 
      n25917, n25918, n25919, n25920, n25921, n25922, n25923, n25924, n25925, 
      n25926, n25927, n25928, n25929, n25930, n25931, n25932, n25933, n25934, 
      n25935, n25936, n25937, n25938, n25939, n25940, n25941, n25942, n25943, 
      n25944, n25945, n25946, n25947, n25948, n25949, n25950, n25951, n25952, 
      n25953, n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961, 
      n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969, n25970, 
      n25971, n25972, n25973, n25974, n25975, n25976, n25977, n25978, n25979, 
      n25980, n25981, n25982, n25983, n25984, n25985, n25986, n25987, n25988, 
      n25989, n25990, n25991, n25992, n25993, n25994, n25995, n25996, n25997, 
      n25998, n25999, n26000, n26001, n26002, n26003, n26004, n26005, n26006, 
      n26007, n26008, n26009, n26010, n26011, n26012, n26013, n26014, n26015, 
      n26016, n26017, n26018, n26019, n26020, n26021, n26022, n26023, n26024, 
      n26025, n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033, 
      n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041, n26042, 
      n26043, n26044, n26045, n26046, n26047, n26048, n26049, n26050, n26051, 
      n26052, n26053, n26054, n26055, n26056, n26057, n26058, n26059, n26060, 
      n26061, n26062, n26063, n26064, n26065, n26066, n26067, n26068, n26069, 
      n26070, n26071, n26072, n26073, n26074, n26075, n26076, n26077, n26078, 
      n26079, n26080, n26081, n26082, n26083, n26084, n26085, n26086, n26087, 
      n26088, n26089, n26090, n26091, n26092, n26093, n26094, n26095, n26096, 
      n26097, n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105, 
      n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113, n26114, 
      n26115, n26116, n26117, n26118, n26119, n26120, n26121, n26122, n26123, 
      n26124, n26125, n26126, n26127, n26128, n26129, n26130, n26131, n26132, 
      n26133, n26134, n26135, n26136, n26137, n26138, n26139, n26140, n26141, 
      n26142, n26143, n26144, n26145, n26146, n26147, n26148, n26149, n26150, 
      n26151, n26152, n26153, n26154, n26155, n26156, n26157, n26158, n26159, 
      n26160, n26161, n26162, n26163, n26164, n26165, n26166, n26167, n26168, 
      n26169, n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177, 
      n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185, n26186, 
      n26187, n26188, n26189, n26190, n26191, n26192, n26193, n26194, n26195, 
      n26196, n26197, n26198, n26199, n26200, n26201, n26202, n26203, n26204, 
      n26205, n26206, n26207, n26208, n26209, n26210, n26211, n26212, n26213, 
      n26214, n26215, n26216, n26217, n26218, n26219, n26220, n26221, n26222, 
      n26223, n26224, n26225, n26226, n26227, n26228, n26229, n26230, n26231, 
      n26232, n26233, n26234, n26235, n26236, n26237, n26238, n26239, n26240, 
      n26241, n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249, 
      n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257, n26258, 
      n26259, n26260, n26261, n26262, n26263, n26264, n26265, n26266, n26267, 
      n26268, n26269, n26270, n26271, n26272, n26273, n26274, n26275, n26276, 
      n26277, n26278, n26279, n26280, n26281, n26282, n26283, n26284, n26285, 
      n26286, n26287, n26288, n26289, n26290, n26291, n26292, n26293, n26294, 
      n26295, n26296, n26297, n26298, n26299, n26300, n26301, n26302, n26303, 
      n26304, n26305, n26306, n26307, n26308, n26309, n26310, n26311, n26312, 
      n26313, n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321, 
      n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329, n26330, 
      n26331, n26332, n26333, n26334, n26335, n26336, n26337, n26338, n26339, 
      n26340, n26341, n26342, n26343, n26344, n26345, n26346, n26347, n26348, 
      n26349, n26350, n26351, n26352, n26353, n26354, n26355, n26356, n26357, 
      n26359, n26361, n26362, n26363, n26364, n26366, n26368, n26369, n26370, 
      n26371, n26373, n26375, n26376, n26377, n26378, n26379, n26380, n26381, 
      n26382, n26383, n26384, n26385, n26386, n26387, n26388, n26389, n26390, 
      n26391, n26392, n26393, n26394, n26397, n26400, n26403, n26404, n26405, 
      n26406, n26407, n26408, n26409, n26410, n26411, n26412, n26413, n26414, 
      n26415, n26416, n26417, n26418, n26419, n26420, n26423, n26426, n26429, 
      n26430, n26431, n26432, n26433, n26434, n26435, n26436, n26437, n26438, 
      n26439, n26440, n26441, n26442, n26443, n26444, n26445, n26446, n26449, 
      n26452, n26455, n26456, n26457, n26458, n26459, n26460, n26461, n26462, 
      n26463, n26464, n26465, n26466, n26467, n26468, n26469, n26470, n26471, 
      n26472, n26475, n26478, n26481, n26482, n26483, n26484, n26485, n26486, 
      n26487, n26488, n26489, n26490, n26491, n26492, n26493, n26494, n26495, 
      n26496, n26497, n26498, n26501, n26504, n26507, n26508, n26509, n26510, 
      n26511, n26512, n26513, n26514, n26515, n26516, n26517, n26518, n26519, 
      n26520, n26521, n26522, n26523, n26524, n26527, n26530, n26533, n26534, 
      n26535, n26536, n26537, n26538, n26539, n26540, n26541, n26542, n26543, 
      n26544, n26545, n26546, n26547, n26548, n26549, n26550, n26553, n26556, 
      n26559, n26560, n26561, n26562, n26563, n26564, n26565, n26566, n26567, 
      n26568, n26569, n26570, n26571, n26572, n26573, n26574, n26575, n26576, 
      n26579, n26582, n26585, n26586, n26587, n26588, n26589, n26590, n26591, 
      n26592, n26593, n26594, n26595, n26596, n26597, n26598, n26599, n26600, 
      n26601, n26602, n26605, n26608, n26611, n26612, n26613, n26614, n26615, 
      n26616, n26617, n26618, n26619, n26620, n26621, n26622, n26623, n26624, 
      n26625, n26626, n26627, n26628, n26631, n26634, n26637, n26638, n26639, 
      n26640, n26641, n26642, n26643, n26644, n26645, n26646, n26647, n26648, 
      n26649, n26650, n26651, n26652, n26653, n26654, n26657, n26660, n26663, 
      n26664, n26665, n26666, n26667, n26668, n26669, n26670, n26671, n26672, 
      n26673, n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26683, 
      n26686, n26689, n26690, n26691, n26692, n26693, n26694, n26695, n26696, 
      n26697, n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705, 
      n26706, n26709, n26712, n26715, n26716, n26717, n26718, n26719, n26720, 
      n26721, n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729, 
      n26730, n26731, n26732, n26735, n26738, n26741, n26742, n26743, n26744, 
      n26745, n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26753, 
      n26754, n26755, n26756, n26757, n26758, n26761, n26764, n26767, n26768, 
      n26769, n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777, 
      n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26787, n26790, 
      n26793, n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801, 
      n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809, n26810, 
      n26813, n26816, n26819, n26820, n26821, n26822, n26823, n26824, n26825, 
      n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833, n26834, 
      n26835, n26836, n26839, n26842, n26845, n26846, n26847, n26848, n26849, 
      n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857, n26858, 
      n26859, n26860, n26861, n26862, n26865, n26868, n26871, n26872, n26873, 
      n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881, n26882, 
      n26883, n26884, n26885, n26886, n26887, n26888, n26891, n26894, n26897, 
      n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905, n26906, 
      n26907, n26908, n26909, n26910, n26911, n26912, n26913, n26914, n26917, 
      n26920, n26923, n26924, n26925, n26926, n26927, n26928, n26929, n26930, 
      n26931, n26932, n26933, n26934, n26935, n26936, n26937, n26938, n26939, 
      n26940, n26943, n26946, n26949, n26950, n26951, n26952, n26953, n26954, 
      n26955, n26956, n26957, n26958, n26959, n26960, n26961, n26962, n26963, 
      n26964, n26965, n26966, n26969, n26972, n26975, n26976, n26977, n26978, 
      n26979, n26980, n26981, n26982, n26983, n26984, n26985, n26986, n26987, 
      n26988, n26989, n26990, n26991, n26992, n26995, n26998, n27001, n27002, 
      n27003, n27004, n27005, n27006, n27007, n27008, n27009, n27010, n27011, 
      n27012, n27013, n27014, n27015, n27016, n27017, n27018, n27021, n27024, 
      n27027, n27028, n27029, n27030, n27031, n27032, n27033, n27034, n27035, 
      n27036, n27037, n27038, n27039, n27040, n27041, n27042, n27043, n27044, 
      n27047, n27050, n27053, n27054, n27055, n27056, n27057, n27058, n27059, 
      n27060, n27061, n27062, n27063, n27064, n27065, n27066, n27067, n27068, 
      n27069, n27070, n27073, n27076, n27079, n27080, n27081, n27082, n27083, 
      n27084, n27085, n27086, n27087, n27088, n27089, n27090, n27091, n27092, 
      n27093, n27094, n27095, n27096, n27099, n27102, n27105, n27106, n27107, 
      n27108, n27109, n27110, n27111, n27112, n27113, n27114, n27115, n27116, 
      n27117, n27118, n27119, n27120, n27121, n27122, n27125, n27128, n27131, 
      n27132, n27133, n27134, n27135, n27136, n27137, n27138, n27139, n27140, 
      n27141, n27142, n27143, n27144, n27145, n27146, n27147, n27148, n27151, 
      n27154, n27157, n27158, n27159, n27160, n27161, n27162, n27163, n27164, 
      n27165, n27166, n27167, n27168, n27169, n27170, n27171, n27172, n27173, 
      n27174, n27177, n27180, n27183, n27184, n27185, n27186, n27187, n27188, 
      n27189, n27190, n27191, n27192, n27193, n27194, n27195, n27196, n27197, 
      n27198, n27199, n27200, n27203, n27206, n27209, n27210, n27211, n27212, 
      n27213, n27214, n27215, n27216, n27217, n27218, n27219, n27220, n27221, 
      n27222, n27223, n27224, n27225, n27226, n27229, n27232, n27235, n27236, 
      n27237, n27238, n27239, n27240, n27241, n27242, n27243, n27244, n27245, 
      n27246, n27247, n27248, n27249, n27250, n27251, n27252, n27255, n27258, 
      n27261, n27262, n27263, n27264, n27265, n27266, n27267, n27268, n27269, 
      n27270, n27271, n27272, n27273, n27274, n27275, n27276, n27277, n27278, 
      n27281, n27284, n27287, n27288, n27289, n27290, n27291, n27292, n27293, 
      n27294, n27295, n27296, n27297, n27298, n27299, n27300, n27301, n27302, 
      n27303, n27304, n27307, n27310, n27313, n27314, n27315, n27316, n27317, 
      n27318, n27319, n27320, n27321, n27322, n27323, n27324, n27325, n27326, 
      n27327, n27328, n27329, n27330, n27333, n27336, n27339, n27340, n27341, 
      n27342, n27343, n27344, n27345, n27346, n27347, n27348, n27349, n27350, 
      n27351, n27352, n27353, n27354, n27355, n27356, n27359, n27362, n27365, 
      n27366, n27367, n27368, n27369, n27370, n27371, n27372, n27373, n27374, 
      n27375, n27376, n27377, n27378, n27379, n27380, n27381, n27382, n27385, 
      n27388, n27391, n27392, n27393, n27394, n27395, n27396, n27397, n27398, 
      n27399, n27400, n27401, n27402, n27403, n27404, n27405, n27406, n27407, 
      n27408, n27411, n27414, n27417, n27418, n27419, n27420, n27421, n27422, 
      n27423, n27424, n27425, n27426, n27427, n27428, n27429, n27430, n27431, 
      n27432, n27433, n27434, n27437, n27440, n27443, n27444, n27445, n27446, 
      n27447, n27448, n27449, n27450, n27451, n27452, n27453, n27454, n27455, 
      n27456, n27457, n27458, n27459, n27460, n27463, n27466, n27469, n27470, 
      n27471, n27472, n27473, n27474, n27475, n27476, n27477, n27478, n27479, 
      n27480, n27481, n27482, n27483, n27484, n27485, n27486, n27489, n27492, 
      n27495, n27496, n27497, n27498, n27499, n27500, n27501, n27502, n27503, 
      n27504, n27505, n27506, n27507, n27508, n27509, n27510, n27511, n27512, 
      n27515, n27518, n27521, n27522, n27523, n27524, n27525, n27526, n27527, 
      n27528, n27529, n27530, n27531, n27532, n27533, n27534, n27535, n27536, 
      n27537, n27538, n27541, n27544, n27547, n27548, n27549, n27550, n27551, 
      n27552, n27553, n27554, n27555, n27556, n27557, n27558, n27559, n27560, 
      n27561, n27562, n27563, n27564, n27567, n27570, n27573, n27574, n27575, 
      n27576, n27577, n27578, n27579, n27580, n27581, n27582, n27583, n27584, 
      n27585, n27586, n27587, n27588, n27589, n27590, n27593, n27596, n27599, 
      n27600, n27601, n27602, n27603, n27604, n27605, n27606, n27607, n27608, 
      n27609, n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27619, 
      n27622, n27625, n27626, n27627, n27628, n27629, n27630, n27631, n27632, 
      n27633, n27634, n27635, n27636, n27637, n27638, n27639, n27640, n27641, 
      n27642, n27645, n27648, n27651, n27652, n27653, n27654, n27655, n27656, 
      n27657, n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665, 
      n27666, n27667, n27668, n27671, n27674, n27677, n27678, n27679, n27680, 
      n27681, n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689, 
      n27690, n27691, n27692, n27693, n27694, n27697, n27700, n27703, n27704, 
      n27705, n27706, n27707, n27708, n27709, n27710, n27711, n27712, n27713, 
      n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27723, n27726, 
      n27729, n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737, 
      n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745, n27746, 
      n27749, n27752, n27755, n27756, n27757, n27758, n27759, n27760, n27761, 
      n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769, n27770, 
      n27771, n27772, n27775, n27778, n27781, n27782, n27783, n27784, n27785, 
      n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793, n27794, 
      n27795, n27796, n27797, n27798, n27801, n27804, n27807, n27808, n27809, 
      n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817, n27818, 
      n27819, n27820, n27821, n27822, n27823, n27824, n27827, n27830, n27833, 
      n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841, n27842, 
      n27843, n27844, n27845, n27846, n27847, n27848, n27849, n27850, n27853, 
      n27856, n27859, n27860, n27861, n27862, n27863, n27864, n27865, n27866, 
      n27867, n27868, n27869, n27870, n27871, n27872, n27873, n27874, n27875, 
      n27876, n27879, n27882, n27885, n27886, n27887, n27888, n27889, n27890, 
      n27891, n27892, n27893, n27894, n27895, n27896, n27897, n27898, n27899, 
      n27900, n27901, n27902, n27905, n27908, n27911, n27912, n27913, n27914, 
      n27915, n27916, n27917, n27918, n27919, n27920, n27921, n27922, n27923, 
      n27924, n27925, n27926, n27927, n27928, n27931, n27934, n27937, n27938, 
      n27939, n27940, n27941, n27942, n27943, n27944, n27945, n27946, n27947, 
      n27948, n27949, n27950, n27951, n27952, n27953, n27954, n27957, n27960, 
      n27963, n27964, n27965, n27966, n27967, n27968, n27969, n27970, n27971, 
      n27972, n27973, n27974, n27975, n27976, n27977, n27978, n27979, n27980, 
      n27983, n27986, n27989, n27990, n27991, n27992, n27993, n27994, n27995, 
      n27996, n27997, n27998, n27999, n28000, n28001, n28002, n28003, n28004, 
      n28005, n28006, n28007, n28008, n28009, n28010, n28011, n28012, n28013, 
      n28014, n28015, n28016, n28017, n28018, n28019, n28020, n28023, n28024, 
      n28027, n28028, n28029, n28032, n28033, n28034, n28035, n28036, n28037, 
      n28038, n28039, n28040, n28041, n28042, n28043, n28044, n28045, n28046, 
      n28047, n28048, n28049, n28050, n28051, n28052, n28053, n28054, n28055, 
      n28056, n28057, n28058, n28059, n28060, n28061, n28062, n28063, n28064, 
      n28065, n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28073, 
      n28074, n28075, n28076, n28077, n28078, n28079, n28080, n28081, n28082, 
      n28083, n28084, n28085, n28086, n28087, n28088, n28089, n28090, n28091, 
      n28092, n28093, n28094, n28095, n28096, n28097, n28098, n28099, n28100, 
      n28101, n28102, n28103, n28104, n28105, n28106, n28107, n28108, n28109, 
      n28110, n28111, n28112, n28113, n28114, n28115, n28116, n28117, n28118, 
      n28119, n28120, n28121, n28122, n28123, n28124, n28125, n28126, n28127, 
      n28128, n28129, n28130, n28131, n28132, n28133, n28134, n28135, n28136, 
      n28137, n28138, n28139, n28140, n28141, n28142, n28143, n28144, n28145, 
      n28146, n28147, n28148, n28149, n28150, n28151, n28152, n28153, n28154, 
      n28155, n28156, n28157, n28158, n28159, n28160, n28161, n28162, n28163, 
      n28164, n28165, n28166, n28167, n28168, n28169, n28170, n28171, n28172, 
      n28173, n28174, n28175, n28176, n28177, n28178, n28179, n28180, n28181, 
      n28182, n28183, n28184, n28185, n28186, n28187, n28188, n28189, n28190, 
      n28191, n28192, n28193, n28194, n28195, n28196, n28197, n28198, n28199, 
      n28200, n28201, n28202, n28203, n28204, n28205, n28206, n28207, n28208, 
      n28209, n28210, n28211, n28212, n28213, n28214, n28215, n28216, n28217, 
      n28218, n28219, n28220, n28221, n28222, n28223, n28224, n28225, n28226, 
      n28227, n28228, n28229, n28230, n28231, n28232, n28233, n28234, n28235, 
      n28236, n28237, n28238, n28239, n28240, n28241, n28242, n28243, n28244, 
      n28245, n28246, n28247, n28248, n28249, n28250, n28251, n28252, n28253, 
      n28254, n28255, n28256, n28257, n28258, n28259, n28260, n28261, n28262, 
      n28263, n28264, n28265, n28266, n28267, n28268, n28269, n28270, n28271, 
      n28272, n28273, n28274, n28275, n28276, n28277, n28278, n28279, n28280, 
      n28281, n28282, n28283, n28284, n28285, n28286, n28287, n28288, n28289, 
      n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297, n28298, 
      n28299, n28300, n28301, n28302, n28303, n28304, n28305, n28306, n28307, 
      n28308, n28309, n28310, n28311, n28312, n28313, n28314, n28315, n28316, 
      n28317, n28318, n28319, n28320, n28321, n28322, n28323, n28324, n28325, 
      n28326, n28327, n28328, n28329, n28330, n28331, n28332, n28333, n28334, 
      n28335, n28336, n28337, n28338, n28339, n28340, n28341, n28342, n28343, 
      n28344, n28345, n28346, n28347, n28348, n28349, n28350, n28351, n28352, 
      n28353, n28354, n28355, n28356, n28357, n28358, n28359, n28360, n28361, 
      n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369, n28370, 
      n28371, n28372, n28373, n28374, n28375, n28376, n28377, n28378, n28379, 
      n28380, n28381, n28382, n28383, n28384, n28385, n28386, n28387, n28388, 
      n28389, n28390, n28391, n28392, n28393, n28394, n28395, n28396, n28397, 
      n28398, n28399, n28400, n28401, n28402, n28403, n28404, n28405, n28406, 
      n28407, n28408, n28409, n28410, n28411, n28412, n28413, n28414, n28415, 
      n28416, n28417, n28418, n28419, n28420, n28421, n28422, n28423, n28424, 
      n28425, n28426, n28427, n28428, n28429, n28430, n28431, n28432, n28433, 
      n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28441, n28442, 
      n28443, n28444, n28445, n28446, n28447, n28448, n28449, n28450, n28451, 
      n28452, n28453, n28454, n28455, n28456, n28457, n28458, n28459, n28460, 
      n28461, n28462, n28463, n28464, n28465, n28466, n28467, n28468, n28469, 
      n28470, n28471, n28472, n28473, n28474, n28475, n28476, n28477, n28478, 
      n28479, n28480, n28481, n28482, n28483, n28484, n28485, n28486, n28487, 
      n28488, n28489, n28490, n28491, n28492, n28493, n28494, n28495, n28496, 
      n28497, n28498, n28499, n28500, n28501, n28502, n28503, n28504, n28505, 
      n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513, n28514, 
      n28515, n28516, n28517, n28518, n28519, n28520, n28521, n28522, n28523, 
      n28524, n28525, n28526, n28527, n28528, n28529, n28530, n28531, n28532, 
      n28533, n28534, n28535, n28536, n28537, n28538, n28539, n28540, n28541, 
      n28542, n28543, n28544, n28545, n28546, n28547, n28548, n28549, n28550, 
      n28551, n28552, n28553, n28554, n28555, n28556, n28557, n28558, n28559, 
      n28560, n28561, n28562, n28563, n28564, n28565, n28566, n28567, n28568, 
      n28569, n28570, n28571, n28572, n28573, n28574, n28575, n28576, n28577, 
      n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585, n28586, 
      n28587, n28588, n28589, n28590, n28591, n28592, n28593, n28594, n28595, 
      n28596, n28597, n28598, n28599, n28600, n28601, n28602, n28603, n28604, 
      n28605, n28606, n28607, n28608, n28609, n28610, n28611, n28612, n28613, 
      n28614, n28615, n28616, n28617, n28618, n28619, n28620, n28621, n28622, 
      n28623, n28624, n28625, n28626, n28627, n28628, n28629, n28630, n28631, 
      n28632, n28633, n28634, n28635, n28636, n28637, n28638, n28639, n28640, 
      n28641, n28642, n28643, n28644, n28645, n28646, n28647, n28648, n28649, 
      n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657, n28658, 
      n28659, n28660, n28661, n28662, n28663, n28664, n28665, n28666, n28667, 
      n28668, n28669, n28670, n28671, n28672, n28673, n28674, n28675, n28676, 
      n28677, n28678, n28679, n28680, n28681, n28682, n28683, n28684, n28685, 
      n28686, n28687, n28688, n28689, n28690, n28691, n28692, n28693, n28694, 
      n28695, n28696, n28697, n28698, n28699, n28700, n28701, n28702, n28703, 
      n28704, n28705, n28706, n28707, n28708, n28709, n28710, n28711, n28712, 
      n28713, n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721, 
      n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729, n28730, 
      n28731, n28732, n28733, n28734, n28735, n28736, n28737, n28738, n28739, 
      n28740, n28741, n28742, n28743, n28744, n28745, n28746, n28747, n28748, 
      n28749, n28750, n28751, n28752, n28753, n28754, n28755, n28756, n28757, 
      n28758, n28759, n28760, n28761, n28762, n28763, n28764, n28765, n28766, 
      n28767, n28768, n28769, n28770, n28771, n28772, n28773, n28774, n28775, 
      n28776, n28777, n28778, n28779, n28780, n28781, n28782, n28783, n28784, 
      n28785, n28786, n28787, n28788, n28789, n28790, n28791, n28792, n28793, 
      n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801, n28802, 
      n28803, n28804, n28805, n28806, n28807, n28808, n28809, n28810, n28811, 
      n28812, n28813, n28814, n28815, n28816, n28817, n28818, n28819, n28820, 
      n28821, n28822, n28823, n28824, n28825, n28826, n28827, n28828, n28829, 
      n28830, n28831, n28832, n28833, n28834, n28835, n28836, n28837, n28838, 
      n28839, n28840, n28841, n28842, n28843, n28844, n28845, n28846, n28847, 
      n28848, n28849, n28850, n28851, n28852, n28853, n28854, n28855, n28856, 
      n28857, n28858, n28859, n28860, n28861, n28862, n28863, n28864, n28865, 
      n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873, n28874, 
      n28875, n28876, n28877, n28878, n28879, n28880, n28881, n28882, n28883, 
      n28884, n28885, n28886, n28887, n28888, n28889, n28890, n28891, n28892, 
      n28893, n28894, n28895, n28896, n28897, n28898, n28899, n28900, n28901, 
      n28902, n28903, n28904, n28905, n28906, n28907, n28908, n28909, n28910, 
      n28911, n28912, n28913, n28914, n28915, n28916, n28917, n28918, n28919, 
      n28920, n28921, n28922, n28923, n28924, n28925, n28926, n28927, n28928, 
      n28929, n28930, n28931, n28932, n28933, n28934, n28935, n28936, n28937, 
      n28938, n28939, n28940, n28941, n28942, n28943, n28944, n28945, n28946, 
      n28947, n28948, n28949, n28950, n28951, n28952, n28953, n28954, n28955, 
      n28956, n28957, n28958, n28959, n28960, n28961, n28962, n28963, n28964, 
      n28965, n28966, n28967, n28968, n28969, n28970, n28971, n28972, n28973, 
      n28974, n28975, n28976, n28977, n28978, n28979, n28980, n28981, n28982, 
      n28983, n28984, n28985, n28986, n28987, n28988, n28989, n28990, n28991, 
      n28992, n28993, n28994, n28995, n28996, n28997, n28998, n28999, n29000, 
      n29001, n29002, n29003, n29004, n29005, n29006, n29007, n29008, n29009, 
      n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017, n29018, 
      n29019, n29020, n29021, n29022, n29023, n29024, n29025, n29026, n29027, 
      n29028, n29029, n29030, n29031, n29032, n29033, n29034, n29035, n29036, 
      n29037, n29038, n29039, n29040, n29041, n29042, n29043, n29044, n29045, 
      n29046, n29047, n29048, n29049, n29050, n29051, n29052, n29053, n29054, 
      n29055, n29056, n29057, n29058, n29059, n29060, n29061, n29062, n29063, 
      n29064, n29065, n29066, n29067, n29068, n29069, n29070, n29071, n29072, 
      n29073, n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081, 
      n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089, n29090, 
      n29091, n29092, n29093, n29094, n29095, n29096, n29097, n29098, n29099, 
      n29100, n29101, n29102, n29103, n29104, n29105, n29106, n29107, n29108, 
      n29109, n29110, n29111, n29112, n29113, n29114, n29115, n29116, n29117, 
      n29118, n29119, n29120, n29121, n29122, n29123, n29124, n29125, n29126, 
      n29127, n29128, n29129, n29130, n29131, n29132, n29133, n29134, n29135, 
      n29136, n29137, n29138, n29139, n29140, n29141, n29142, n29143, n29144, 
      n29145, n29146, n29147, n29148, n29149, n29150, n29151, n29152, n29153, 
      n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161, n29162, 
      n29163, n29164, n29165, n29166, n29167, n29168, n29169, n29170, n29171, 
      n29172, n29173, n29174, n29175, n29176, n29177, n29178, n29179, n29180, 
      n29181, n29182, n29183, n29184, n29185, n29186, n29187, n29188, n29189, 
      n29190, n29191, n29192, n29193, n29194, n29195, n29196, n29197, n29198, 
      n29199, n29200, n29201, n29202, n29203, n29204, n29205, n29206, n29207, 
      n29208, n29209, n29210, n29211, n29212, n29213, n29214, n29215, n29216, 
      n29217, n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29225, 
      n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233, n29234, 
      n29235, n29236, n29237, n29238, n29239, n29240, n29241, n29242, n29243, 
      n29244, n29245, n29246, n29247, n29248, n29249, n29250, n29251, n29252, 
      n29253, n29254, n29255, n29256, n29257, n29258, n29259, n29260, n29261, 
      n29262, n29263, n29264, n29265, n29266, n29267, n29268, n29269, n29270, 
      n29271, n29272, n29273, n29274, n29275, n29276, n29277, n29278, n29279, 
      n29280, n29281, n29282, n29283, n29284, n29285, n29286, n29287, n29288, 
      n29289, n29290, n29291, n29292, n29293, n29294, n29295, n29296, n29297, 
      n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305, n29306, 
      n29307, n29308, n29309, n29310, n29311, n29312, n29313, n29314, n29315, 
      n29316, n29317, n29318, n29319, n29320, n29321, n29322, n29323, n29324, 
      n29325, n29326, n29327, n29328, n29329, n29330, n29331, n29332, n29333, 
      n29334, n29335, n29336, n29337, n29338, n29339, n29340, n29341, n29342, 
      n29343, n29344, n29345, n29346, n29347, n29348, n29349, n29350, n29351, 
      n29352, n29353, n29354, n29355, n29356, n29357, n29358, n29359, n29360, 
      n29361, n29362, n29363, n29364, n29365, n29366, n29367, n29368, n29369, 
      n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377, n29378, 
      n29379, n29380, n29381, n29382, n29383, n29384, n29385, n29386, n29387, 
      n29388, n29389, n29390, n29391, n29392, n29393, n29394, n29395, n29396, 
      n29397, n29398, n29399, n29400, n29401, n29402, n29403, n29404, n29405, 
      n29406, n29407, n29408, n29409, n29410, n29411, n29412, n29413, n29414, 
      n29415, n29416, n29417, n29418, n29419, n29420, n29421, n29422, n29423, 
      n29424, n29425, n29426, n29427, n29428, n29429, n29430, n29431, n29432, 
      n29433, n29434, n29435, n29436, n29437, n29438, n29439, n29440, n29441, 
      n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449, n29450, 
      n29451, n29452, n29453, n29454, n29455, n29456, n29457, n29458, n29459, 
      n29460, n29461, n29462, n29463, n29464, n29465, n29466, n29467, n29468, 
      n29469, n29470, n29471, n29472, n29473, n29474, n29475, n29476, n29477, 
      n29478, n29479, n29480, n29481, n29482, n29483, n29484, n29485, n29486, 
      n29487, n29488, n29489, n29490, n29491, n29492, n29493, n29494, n29495, 
      n29496, n29497, n29498, n29499, n29500, n29501, n29502, n29503, n29504, 
      n29505, n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513, 
      n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521, n29522, 
      n29523, n29524, n29525, n29526, n29527, n29528, n29529, n29530, n29531, 
      n29532, n29533, n29534, n29535, n29536, n29537, n29538, n29539, n29540, 
      n29541, n29542, n29543, n29544, n29545, n29546, n29547, n29548, n29549, 
      n29550, n29551, n29552, n29553, n29554, n29555, n29556, n29557, n29558, 
      n29559, n29560, n29561, n29562, n29563, n29564, n29565, n29566, n29567, 
      n29568, n29569, n29570, n29571, n29572, n29573, n29574, n29575, n29576, 
      n29577, n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585, 
      n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593, n29594, 
      n29595, n29596, n29597, n29598, n29599, n29600, n29601, n29602, n29603, 
      n29604, n29605, n29606, n29607, n29608, n29609, n29610, n29611, n29612, 
      n29613, n29614, n29615, n29616, n29617, n29618, n29619, n29620, n29621, 
      n29622, n29623, n29624, n29625, n29626, n29627, n29628, n29629, n29630, 
      n29631, n29632, n29633, n29634, n29635, n29636, n29637, n29638, n29639, 
      n29640, n29641, n29642, n29643, n29644, n29645, n29646, n29647, n29648, 
      n29649, n29650, n29651, n29652, n29653, n29654, n29655, n29656, n29657, 
      n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665, n29666, 
      n29667, n29668, n29669, n29670, n29671, n29672, n29673, n29674, n29675, 
      n29676, n29677, n29678, n29679, n29680, n29681, n29682, n29683, n29684, 
      n29685, n29686, n29687, n29688, n29689, n29690, n29691, n29692, n29693, 
      n29694, n29695, n29696, n29697, n29698, n29699, n29700, n29701, n29702, 
      n29703, n29704, n29705, n29706, n29707, n29708, n29709, n29710, n29711, 
      n29712, n29713, n29714, n29715, n29716, n29717, n29718, n29719, n29720, 
      n29721, n29722, n29723, n29724, n29725, n29726, n29727, n29728, n29729, 
      n29730, n29731, n29732, n29733, n29734, n29735, n29736, n29737, n29738, 
      n29739, n29740, n29741, n29742, n29743, n29744, n29745, n29746, n29747, 
      n29748, n29749, n29750, n29751, n29752, n29753, n29754, n29755, n29756, 
      n29757, n29758, n29759, n29760, n29761, n29762, n29763, n29764, n29765, 
      n29766, n29767, n29768, n29769, n29770, n29771, n29772, n29773, n29774, 
      n29775, n29776, n29777, n29778, n29779, n29780, n29781, n29782, n29783, 
      n29784, n29785, n29786, n29787, n29788, n29789, n29790, n29791, n29792, 
      n29793, n29794, n29795, n29796, n29797, n29798, n29799, n29800, n29801, 
      n29802, n29803, n29804, n29805, n29806, n29807, n29808, n29809, n29810, 
      n29811, n29812, n29813, n29814, n29815, n29816, n29817, n29818, n29819, 
      n29820, n29821, n29822, n29823, n29824, n29825, n29826, n29827, n29828, 
      n29829, n29830, n29831, n29832, n29833, n29834, n29835, n29836, n29837, 
      n29838, n29839, n29840, n29841, n29842, n29843, n29844, n29845, n29846, 
      n29847, n29848, n29849, n29850, n29851, n29852, n29853, n29854, n29855, 
      n29856, n29857, n29858, n29859, n29860, n29861, n29862, n29863, n29864, 
      n29865, n29866, n29867, n29868, n29869, n29870, n29871, n29872, n29873, 
      n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881, n29882, 
      n29883, n29884, n29885, n29886, n29887, n29888, n29889, n29890, n29891, 
      n29892, n29893, n29894, n29895, n29896, n29897, n29898, n29899, n29900, 
      n29901, n29902, n29903, n29904, n29905, n29906, n29907, n29908, n29909, 
      n29910, n29911, n29912, n29913, n29914, n29915, n29916, n29917, n29918, 
      n29919, n29920, n29921, n29922, n29923, n29924, n29925, n29926, n29927, 
      n29928, n29929, n29930, n29931, n29932, n29933, n29934, n29935, n29936, 
      n29937, n29938, n29939, n29940, n29941, n29942, n29943, n29944, n29945, 
      n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953, n29954, 
      n29955, n29956, n29957, n29958, n29959, n29960, n29961, n29962, n29963, 
      n29964, n29965, n29966, n29967, n29968, n29969, n29970, n29971, n29972, 
      n29973, n29974, n29975, n29976, n29977, n29978, n29979, n29980, n29981, 
      n29982, n29983, n29984, n29985, n29986, n29987, n29988, n29989, n29990, 
      n29991, n29992, n29993, n29994, n29995, n29996, n29997, n29998, n29999, 
      n30000, n30001, n30002, n30003, n30004, n30005, n30006, n30007, n30008, 
      n30009, n30010, n30011, n30012, n30013, n30014, n30015, n30016, n30017, 
      n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025, n30026, 
      n30027, n30028, n30029, n30030, n30031, n30032, n30033, n30034, n30035, 
      n30036, n30037, n30038, n30039, n30040, n30041, n30042, n30043, n30044, 
      n30045, n30046, n30047, n30048, n30049, n30050, n30051, n30052, n30053, 
      n30054, n30055, n30056, n30057, n30058, n30059, n30060, n30061, n30062, 
      n30063, n30064, n30065, n30066, n30067, n30068, n30069, n30070, n30071, 
      n30072, n30073, n30074, n30075, n30076, n30077, n30078, n30079, n30080, 
      n30081, n30082, n30083, n30084, n30085, n30086, n30087, n30088, n30089, 
      n30090, n30091, n30092, n30093, n30094, n30095, n30096, n30097, n30098, 
      n30099, n30100, n30101, n30102, n30103, n30104, n30105, n30106, n30107, 
      n30108, n30109, n30110, n30111, n30112, n30113, n30114, n30115, n30116, 
      n30117, n30118, n30119, n30120, n30121, n30122, n30123, n30124, n30125, 
      n30126, n30127, n30128, n30129, n30130, n30131, n30132, n30133, n30134, 
      n30135, n30136, n30137, n30138, n30139, n30140, n30141, n30142, n30143, 
      n30144, n30145, n30146, n30147, n30148, n30149, n30150, n30151, n30152, 
      n30153, n30154, n30155, n30156, n30157, n30158, n30159, n30160, n30161, 
      n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169, n30170, 
      n30171, n30172, n30173, n30174, n30175, n30176, n30177, n30178, n30179, 
      n30180, n30181, n30182, n30183, n30184, n30185, n30186, n30187, n30188, 
      n30189, n30190, n30191, n30192, n30193, n30194, n30195, n30196, n30197, 
      n30198, n30199, n30200, n30201, n30202, n30203, n30204, n30205, n30206, 
      n30207, n30208, n30209, n30210, n30211, n30212, n30213, n30214, n30215, 
      n30216, n30217, n30218, n30219, n30220, n30221, n30222, n30223, n30224, 
      n30225, n30226, n30227, n30228, n30229, n30230, n30231, n30232, n30233, 
      n30234, n30235, n30236, n30237, n30238, n30239, n30240, n30241, n30242, 
      n30243, n30244, n30245, n30246, n30247, n30248, n30249, n30250, n30251, 
      n30252, n30253, n30254, n30255, n30256, n30257, n30258, n30259, n30260, 
      n30261, n30262, n30263, n30264, n30265, n30266, n30267, n30268, n30269, 
      n30270, n30271, n30272, n30273, n30274, n30275, n30276, n30277, n30278, 
      n30279, n30280, n30281, n30282, n30283, n30284, n30285, n30286, n30287, 
      n30288, n30289, n30290, n30291, n30292, n30293, n30294, n30295, n30296, 
      n30297, n30298, n30299, n30300, n30301, n30302, n30303, n30304, n30305, 
      n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313, n30314, 
      n30315, n30316, n30317, n30318, n30319, n30320, n30321, n30322, n30323, 
      n30324, n30325, n30326, n30327, n30328, n30329, n30330, n30331, n30332, 
      n30333, n30334, n30335, n30336, n30337, n30338, n30339, n30340, n30341, 
      n30342, n30343, n30344, n30345, n30346, n30347, n30348, n30349, n30350, 
      n30351, n30352, n30353, n30354, n30355, n30356, n30357, n30358, n30359, 
      n30360, n30361, n30362, n30363, n30364, n30365, n30366, n30367, n30368, 
      n30369, n30370, n30371, n30372, n30373, n30374, n30375, n30376, n30377, 
      n30378, n30379, n30380, n30381, n30382, n30383, n30384, n30385, n30386, 
      n30387, n30388, n30389, n30390, n30391, n30392, n30393, n30394, n30395, 
      n30396, n30397, n30398, n30399, n30400, n30401, n30402, n30403, n30404, 
      n30405, n30406, n30407, n30408, n30409, n30410, n30411, n30412, n30413, 
      n30414, n30415, n30416, n30417, n30418, n30419, n30420, n30421, n30422, 
      n30423, n30424, n30425, n30426, n30427, n30428, n30429, n30430, n30431, 
      n30432, n30433, n30434, n30435, n30436, n30437, n30438, n30439, n30440, 
      n30441, n30442, n30443, n30444, n30445, n30446, n30447, n30448, n30449, 
      n30450, n30451, n30452, n30453, n30454, n30455, n30456, n30457, n30458, 
      n30459, n30460, n30461, n30462, n30463, n30464, n30465, n30466, n30467, 
      n30468, n30469, n30470, n30471, n30472, n30473, n30474, n30475, n30476, 
      n30477, n30478, n30479, n30480, n30481, n30482, n30483, n30484, n30485, 
      n30486, n30487, n30488, n30489, n30490, n30491, n30492, n30493, n30494, 
      n30495, n30496, n30497, n30498, n30499, n30500, n30501, n30502, n30503, 
      n30504, n30505, n30506, n30507, n30508, n30509, n30510, n30511, n30512, 
      n30513, n30514, n30515, n30516, n30517, n30518, n30519, n30520, n30521, 
      n30522, n30523, n30524, n30525, n30526, n30527, n30528, n30529, n30530, 
      n30531, n30532, n30533, n30534, n30535, n30536, n30537, n30538, n30539, 
      n30540, n30541, n30542, n30543, n30544, n30545, n30546, n30547, n30548, 
      n30549, n30550, n30551, n30552, n30553, n30554, n30555, n30556, n30557, 
      n30558, n30559, n30560, n30561, n30562, n30563, n30564, n30565, n30566, 
      n30567, n30568, n30569, n30570, n30571, n30572, n30573, n30574, n30575, 
      n30576, n30577, n30578, n30579, n30580, n30581, n30582, n30583, n30584, 
      n30585, n30586, n30587, n30588, n30589, n30590, n30591, n30592, n30593, 
      n30594, n30595, n30596, n30597, n30598, n30599, n30600, n30601, n30602, 
      n30603, n30604, n30605, n30606, n30607, n30608, n30609, n30610, n30611, 
      n30612, n30613, n30614, n30615, n30616, n30617, n30618, n30619, n30620, 
      n30621, n30622, n30623, n30624, n30625, n30626, n30627, n30628, n30629, 
      n30630, n30631, n30632, n30633, n30634, n30635, n30636, n30637, n30638, 
      n30639, n30640, n30641, n30642, n30643, n30644, n30645, n30646, n30647, 
      n30648, n30649, n30650, n30651, n30652, n30653, n30654, n30655, n30656, 
      n30657, n30658, n30659, n30660, n30661, n30662, n30663, n30664, n30665, 
      n30666, n30667, n30668, n30669, n30670, n30671, n30672, n30673, n30674, 
      n30675, n30676, n30677, n30678, n30679, n30680, n30681, n30682, n30683, 
      n30684, n30685, n30686, n30687, n30688, n30689, n30690, n30691, n30692, 
      n30693, n30694, n30695, n30696, n30697, n30698, n30699, n30700, n30701, 
      n30702, n30703, n30704, n30705, n30706, n30707, n30708, n30709, n30710, 
      n30711, n30712, n30713, n30714, n30715, n30716, n30717, n30718, n30719, 
      n30720, n30721, n30722, n30723, n30724, n30725, n30726, n30727, n30728, 
      n30729, n30730, n30731, n30732, n30733, n30734, n30735, n30736, n30737, 
      n30738, n30739, n30740, n30741, n30742, n30743, n30744, n30745, n30746, 
      n30747, n30748, n30749, n30750, n30751, n30752, n30753, n30754, n30755, 
      n30756, n30757, n30758, n30759, n30760, n30761, n30762, n30763, n30764, 
      n30765, n30766, n30767, n30768, n30769, n30770, n30771, n30772, n30773, 
      n30774, n30775, n30776, n30777, n30778, n30779, n30780, n30781, n30782, 
      n30783, n30784, n30785, n30786, n30787, n30788, n30789, n30790, n30791, 
      n30792, n30793, n30794, n30795, n30796, n30797, n30798, n30799, n30800, 
      n30801, n30802, n30803, n30804, n30805, n30806, n30807, n30808, n30809, 
      n30810, n30811, n30812, n30813, n30814, n30815, n30816, n30817, n30818, 
      n30819, n30820, n30821, n30822, n30823, n30824, n30825, n30826, n30827, 
      n30828, n30829, n30830, n30831, n30832, n30833, n30834, n30835, n30836, 
      n30837, n30838, n30839, n30840, n30841, n30842, n30843, n30844, n30845, 
      n30846, n30847, n30848, n30849, n30850, n30851, n30852, n30853, n30854, 
      n30855, n30856, n30857, n30858, n30859, n30860, n30861, n30862, n30863, 
      n30864, n30865, n30866, n30867, n30868, n30869, n30870, n30871, n30872, 
      n30873, n30874, n30875, n30876, n30877, n30878, n30879, n30880, n30881, 
      n30882, n30883, n30884, n30885, n30886, n30887, n30888, n30889, n30890, 
      n30891, n30892, n30893, n30894, n30895, n30896, n30897, n30898, n30899, 
      n30900, n30901, n30902, n30903, n30904, n30905, n30906, n30907, n30908, 
      n30909, n30910, n30911, n30912, n30913, n30914, n30915, n30916, n30917, 
      n30918, n30919, n30920, n30921, n30922, n30923, n30924, n30925, n30926, 
      n30927, n30928, n30929, n30930, n30931, n30932, n30933, n30934, n30935, 
      n30936, n30937, n30938, n30939, n30940, n30941, n30942, n30943, n30944, 
      n30945, n30946, n30947, n30948, n30949, n30950, n30951, n30952, n30953, 
      n30954, n30955, n30956, n30957, n30958, n30959, n30960, n30961, n30962, 
      n30963, n30964, n30965, n30966, n30967, n30968, n30969, n30970, n30971, 
      n30972, n30973, n30974, n30975, n30976, n30977, n30978, n30979, n30980, 
      n30981, n30982, n30983, n30984, n30985, n30986, n30987, n30988, n30989, 
      n30990, n30991, n30992, n30993, n30994, n30995, n30996, n30997, n30998, 
      n30999, n31000, n31001, n31002, n31003, n31004, n31005, n31006, n31007, 
      n31008, n31009, n31010, n31011, n31012, n31013, n31014, n31015, n31016, 
      n31017, n31018, n31019, n31020, n31021, n31022, n31023, n31024, n31025, 
      n31026, n31027, n31028, n31029, n31030, n31031, n31032, n31033, n31034, 
      n31035, n31036, n31037, n31038, n31039, n31040, n31041, n31042, n31043, 
      n31044, n31045, n31046, n31047, n31048, n31049, n31050, n31051, n31052, 
      n31053, n31054, n31055, n31056, n31057, n31058, n31059, n31060, n31061, 
      n31062, n31063, n31064, n31065, n31066, n31067, n31068, n31069, n31070, 
      n31071, n31072, n31073, n31074, n31075, n31076, n31077, n31078, n31079, 
      n31080, n31081, n31082, n31083, n31084, n31085, n31086, n31087, n31088, 
      n31089, n31090, n31091, n31092, n31093, n31094, n31095, n31096, n31097, 
      n31098, n31099, n31100, n31101, n31102, n31103, n31104, n31105, n31106, 
      n31107, n31108, n31109, n31110, n31111, n31112, n31113, n31114, n31115, 
      n31116, n31117, n31118, n31119, n31120, n31121, n31122, n31123, n31124, 
      n31125, n31126, n31127, n31128, n31129, n31130, n31131, n31132, n31133, 
      n31134, n31135, n31136, n31137, n31138, n31139, n31140, n31141, n31142, 
      n31143, n31144, n31145, n31146, n31147, n31148, n31149, n31150, n31151, 
      n31152, n31153, n31154, n31155, n31156, n31157, n31158, n31159, n31160, 
      n31161, n31162, n31163, n31164, n31165, n31166, n31167, n31168, n31169, 
      n31170, n31171, n31172, n31173, n31174, n31175, n31176, n31177, n31178, 
      n31179, n31180, n31181, n31182, n31183, n31184, n31185, n31186, n31187 : 
      std_logic;

begin
   
   OUT2_tri_enable_reg_63_inst : DFF_X1 port map( D => n7944, CK => CLK, Q => 
                           n5130, QN => n10889);
   OUT2_tri_enable_reg_62_inst : DFF_X1 port map( D => n7943, CK => CLK, Q => 
                           n5132, QN => n10890);
   OUT2_tri_enable_reg_61_inst : DFF_X1 port map( D => n7942, CK => CLK, Q => 
                           n5134, QN => n10891);
   OUT2_tri_enable_reg_60_inst : DFF_X1 port map( D => n7941, CK => CLK, Q => 
                           n5136, QN => n10892);
   OUT2_tri_enable_reg_59_inst : DFF_X1 port map( D => n7940, CK => CLK, Q => 
                           n5138, QN => n10893);
   OUT2_tri_enable_reg_58_inst : DFF_X1 port map( D => n7939, CK => CLK, Q => 
                           n5140, QN => n10894);
   OUT2_tri_enable_reg_57_inst : DFF_X1 port map( D => n7938, CK => CLK, Q => 
                           n5142, QN => n10895);
   OUT2_tri_enable_reg_56_inst : DFF_X1 port map( D => n7937, CK => CLK, Q => 
                           n5144, QN => n10896);
   OUT2_tri_enable_reg_55_inst : DFF_X1 port map( D => n7936, CK => CLK, Q => 
                           n5146, QN => n10897);
   OUT2_tri_enable_reg_54_inst : DFF_X1 port map( D => n7935, CK => CLK, Q => 
                           n5148, QN => n10898);
   OUT2_tri_enable_reg_53_inst : DFF_X1 port map( D => n7934, CK => CLK, Q => 
                           n5150, QN => n10899);
   OUT2_tri_enable_reg_52_inst : DFF_X1 port map( D => n7933, CK => CLK, Q => 
                           n5152, QN => n10900);
   OUT2_tri_enable_reg_51_inst : DFF_X1 port map( D => n7932, CK => CLK, Q => 
                           n5154, QN => n10901);
   OUT2_tri_enable_reg_50_inst : DFF_X1 port map( D => n7931, CK => CLK, Q => 
                           n5156, QN => n10902);
   OUT2_tri_enable_reg_49_inst : DFF_X1 port map( D => n7930, CK => CLK, Q => 
                           n5158, QN => n10903);
   OUT2_tri_enable_reg_48_inst : DFF_X1 port map( D => n7929, CK => CLK, Q => 
                           n5160, QN => n10904);
   OUT2_tri_enable_reg_47_inst : DFF_X1 port map( D => n7928, CK => CLK, Q => 
                           n5162, QN => n10905);
   OUT2_tri_enable_reg_46_inst : DFF_X1 port map( D => n7927, CK => CLK, Q => 
                           n5164, QN => n10906);
   OUT2_tri_enable_reg_45_inst : DFF_X1 port map( D => n7926, CK => CLK, Q => 
                           n5166, QN => n10907);
   OUT2_tri_enable_reg_44_inst : DFF_X1 port map( D => n7925, CK => CLK, Q => 
                           n5168, QN => n10908);
   OUT2_tri_enable_reg_43_inst : DFF_X1 port map( D => n7924, CK => CLK, Q => 
                           n5170, QN => n10909);
   OUT2_tri_enable_reg_42_inst : DFF_X1 port map( D => n7923, CK => CLK, Q => 
                           n5172, QN => n10910);
   OUT2_tri_enable_reg_41_inst : DFF_X1 port map( D => n7922, CK => CLK, Q => 
                           n5174, QN => n10911);
   OUT2_tri_enable_reg_40_inst : DFF_X1 port map( D => n7921, CK => CLK, Q => 
                           n5176, QN => n10912);
   OUT2_tri_enable_reg_39_inst : DFF_X1 port map( D => n7920, CK => CLK, Q => 
                           n5178, QN => n10913);
   OUT2_tri_enable_reg_38_inst : DFF_X1 port map( D => n7919, CK => CLK, Q => 
                           n5180, QN => n10914);
   OUT2_tri_enable_reg_37_inst : DFF_X1 port map( D => n7918, CK => CLK, Q => 
                           n5182, QN => n10915);
   OUT2_tri_enable_reg_36_inst : DFF_X1 port map( D => n7917, CK => CLK, Q => 
                           n5184, QN => n10916);
   OUT2_tri_enable_reg_35_inst : DFF_X1 port map( D => n7916, CK => CLK, Q => 
                           n5186, QN => n10917);
   OUT2_tri_enable_reg_34_inst : DFF_X1 port map( D => n7915, CK => CLK, Q => 
                           n5188, QN => n10918);
   OUT2_tri_enable_reg_33_inst : DFF_X1 port map( D => n7914, CK => CLK, Q => 
                           n5190, QN => n10919);
   OUT2_tri_enable_reg_32_inst : DFF_X1 port map( D => n7913, CK => CLK, Q => 
                           n5192, QN => n10920);
   OUT2_tri_enable_reg_31_inst : DFF_X1 port map( D => n7912, CK => CLK, Q => 
                           n5194, QN => n10921);
   OUT2_tri_enable_reg_30_inst : DFF_X1 port map( D => n7911, CK => CLK, Q => 
                           n5196, QN => n10922);
   OUT2_tri_enable_reg_29_inst : DFF_X1 port map( D => n7910, CK => CLK, Q => 
                           n5198, QN => n10923);
   OUT2_tri_enable_reg_28_inst : DFF_X1 port map( D => n7909, CK => CLK, Q => 
                           n5200, QN => n10924);
   OUT2_tri_enable_reg_27_inst : DFF_X1 port map( D => n7908, CK => CLK, Q => 
                           n5202, QN => n10925);
   OUT2_tri_enable_reg_26_inst : DFF_X1 port map( D => n7907, CK => CLK, Q => 
                           n5204, QN => n10926);
   OUT2_tri_enable_reg_25_inst : DFF_X1 port map( D => n7906, CK => CLK, Q => 
                           n5206, QN => n10927);
   OUT2_tri_enable_reg_24_inst : DFF_X1 port map( D => n7905, CK => CLK, Q => 
                           n5208, QN => n10928);
   OUT2_tri_enable_reg_23_inst : DFF_X1 port map( D => n7904, CK => CLK, Q => 
                           n5210, QN => n10929);
   OUT2_tri_enable_reg_22_inst : DFF_X1 port map( D => n7903, CK => CLK, Q => 
                           n5212, QN => n10930);
   OUT2_tri_enable_reg_21_inst : DFF_X1 port map( D => n7902, CK => CLK, Q => 
                           n5214, QN => n10931);
   OUT2_tri_enable_reg_20_inst : DFF_X1 port map( D => n7901, CK => CLK, Q => 
                           n5216, QN => n10932);
   OUT2_tri_enable_reg_19_inst : DFF_X1 port map( D => n7900, CK => CLK, Q => 
                           n5218, QN => n10933);
   OUT2_tri_enable_reg_18_inst : DFF_X1 port map( D => n7899, CK => CLK, Q => 
                           n5220, QN => n10934);
   OUT2_tri_enable_reg_17_inst : DFF_X1 port map( D => n7898, CK => CLK, Q => 
                           n5222, QN => n10935);
   OUT2_tri_enable_reg_16_inst : DFF_X1 port map( D => n7897, CK => CLK, Q => 
                           n5224, QN => n10936);
   OUT2_tri_enable_reg_15_inst : DFF_X1 port map( D => n7896, CK => CLK, Q => 
                           n5226, QN => n10937);
   OUT2_tri_enable_reg_14_inst : DFF_X1 port map( D => n7895, CK => CLK, Q => 
                           n5228, QN => n10938);
   OUT2_tri_enable_reg_13_inst : DFF_X1 port map( D => n7894, CK => CLK, Q => 
                           n5230, QN => n10939);
   OUT2_tri_enable_reg_12_inst : DFF_X1 port map( D => n7893, CK => CLK, Q => 
                           n5232, QN => n10940);
   OUT2_tri_enable_reg_11_inst : DFF_X1 port map( D => n7892, CK => CLK, Q => 
                           n5234, QN => n10941);
   OUT2_tri_enable_reg_10_inst : DFF_X1 port map( D => n7891, CK => CLK, Q => 
                           n5236, QN => n10942);
   OUT2_tri_enable_reg_9_inst : DFF_X1 port map( D => n7890, CK => CLK, Q => 
                           n5238, QN => n10943);
   OUT2_tri_enable_reg_8_inst : DFF_X1 port map( D => n7889, CK => CLK, Q => 
                           n5240, QN => n10944);
   OUT2_tri_enable_reg_7_inst : DFF_X1 port map( D => n7888, CK => CLK, Q => 
                           n5242, QN => n10945);
   OUT2_tri_enable_reg_6_inst : DFF_X1 port map( D => n7887, CK => CLK, Q => 
                           n5244, QN => n10946);
   OUT2_tri_enable_reg_5_inst : DFF_X1 port map( D => n7886, CK => CLK, Q => 
                           n5246, QN => n10947);
   OUT2_tri_enable_reg_4_inst : DFF_X1 port map( D => n7885, CK => CLK, Q => 
                           n5248, QN => n10948);
   OUT2_tri_enable_reg_3_inst : DFF_X1 port map( D => n7884, CK => CLK, Q => 
                           n5250, QN => n10949);
   OUT2_tri_enable_reg_2_inst : DFF_X1 port map( D => n7883, CK => CLK, Q => 
                           n5252, QN => n10950);
   OUT2_tri_enable_reg_1_inst : DFF_X1 port map( D => n7882, CK => CLK, Q => 
                           n5254, QN => n10951);
   OUT2_tri_enable_reg_0_inst : DFF_X1 port map( D => n7881, CK => CLK, Q => 
                           n5256, QN => n10952);
   REGISTERS_reg_0_63_inst : DFF_X1 port map( D => n7880, CK => CLK, Q => 
                           n15828, QN => n9737);
   REGISTERS_reg_0_62_inst : DFF_X1 port map( D => n7879, CK => CLK, Q => 
                           n15827, QN => n9742);
   REGISTERS_reg_0_61_inst : DFF_X1 port map( D => n7878, CK => CLK, Q => 
                           n15826, QN => n9747);
   REGISTERS_reg_0_60_inst : DFF_X1 port map( D => n7877, CK => CLK, Q => 
                           n15825, QN => n9752);
   REGISTERS_reg_0_59_inst : DFF_X1 port map( D => n7876, CK => CLK, Q => 
                           n15824, QN => n9757);
   REGISTERS_reg_0_58_inst : DFF_X1 port map( D => n7875, CK => CLK, Q => 
                           n15823, QN => n9762);
   REGISTERS_reg_0_57_inst : DFF_X1 port map( D => n7874, CK => CLK, Q => 
                           n15822, QN => n9767);
   REGISTERS_reg_0_56_inst : DFF_X1 port map( D => n7873, CK => CLK, Q => 
                           n15821, QN => n9772);
   REGISTERS_reg_0_55_inst : DFF_X1 port map( D => n7872, CK => CLK, Q => 
                           n15820, QN => n9777);
   REGISTERS_reg_0_54_inst : DFF_X1 port map( D => n7871, CK => CLK, Q => 
                           n15819, QN => n9782);
   REGISTERS_reg_0_53_inst : DFF_X1 port map( D => n7870, CK => CLK, Q => 
                           n15818, QN => n9787);
   REGISTERS_reg_0_52_inst : DFF_X1 port map( D => n7869, CK => CLK, Q => 
                           n15817, QN => n9792);
   REGISTERS_reg_0_51_inst : DFF_X1 port map( D => n7868, CK => CLK, Q => 
                           n15816, QN => n9797);
   REGISTERS_reg_0_50_inst : DFF_X1 port map( D => n7867, CK => CLK, Q => 
                           n15815, QN => n9802);
   REGISTERS_reg_0_49_inst : DFF_X1 port map( D => n7866, CK => CLK, Q => 
                           n15814, QN => n9807);
   REGISTERS_reg_0_48_inst : DFF_X1 port map( D => n7865, CK => CLK, Q => 
                           n15813, QN => n9812);
   REGISTERS_reg_0_47_inst : DFF_X1 port map( D => n7864, CK => CLK, Q => 
                           n15812, QN => n9817);
   REGISTERS_reg_0_46_inst : DFF_X1 port map( D => n7863, CK => CLK, Q => 
                           n15811, QN => n9822);
   REGISTERS_reg_0_45_inst : DFF_X1 port map( D => n7862, CK => CLK, Q => 
                           n15810, QN => n9827);
   REGISTERS_reg_0_44_inst : DFF_X1 port map( D => n7861, CK => CLK, Q => 
                           n15809, QN => n9832);
   REGISTERS_reg_0_43_inst : DFF_X1 port map( D => n7860, CK => CLK, Q => 
                           n15808, QN => n9837);
   REGISTERS_reg_0_42_inst : DFF_X1 port map( D => n7859, CK => CLK, Q => 
                           n15807, QN => n9842);
   REGISTERS_reg_0_41_inst : DFF_X1 port map( D => n7858, CK => CLK, Q => 
                           n15806, QN => n9847);
   REGISTERS_reg_0_40_inst : DFF_X1 port map( D => n7857, CK => CLK, Q => 
                           n15805, QN => n9852);
   REGISTERS_reg_0_39_inst : DFF_X1 port map( D => n7856, CK => CLK, Q => 
                           n15804, QN => n9857);
   REGISTERS_reg_0_38_inst : DFF_X1 port map( D => n7855, CK => CLK, Q => 
                           n15803, QN => n9862);
   REGISTERS_reg_0_37_inst : DFF_X1 port map( D => n7854, CK => CLK, Q => 
                           n15802, QN => n9867);
   REGISTERS_reg_0_36_inst : DFF_X1 port map( D => n7853, CK => CLK, Q => 
                           n15801, QN => n9872);
   REGISTERS_reg_0_35_inst : DFF_X1 port map( D => n7852, CK => CLK, Q => 
                           n15800, QN => n9877);
   REGISTERS_reg_0_34_inst : DFF_X1 port map( D => n7851, CK => CLK, Q => 
                           n15799, QN => n9882);
   REGISTERS_reg_0_33_inst : DFF_X1 port map( D => n7850, CK => CLK, Q => 
                           n15798, QN => n9887);
   REGISTERS_reg_0_32_inst : DFF_X1 port map( D => n7849, CK => CLK, Q => 
                           n15797, QN => n9892);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n7848, CK => CLK, Q => 
                           n15796, QN => n9897);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n7847, CK => CLK, Q => 
                           n15795, QN => n9902);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n7846, CK => CLK, Q => 
                           n15794, QN => n9907);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n7845, CK => CLK, Q => 
                           n15793, QN => n9912);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n7844, CK => CLK, Q => 
                           n15792, QN => n9917);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n7843, CK => CLK, Q => 
                           n15791, QN => n9922);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n7842, CK => CLK, Q => 
                           n15790, QN => n9927);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n7841, CK => CLK, Q => 
                           n15789, QN => n9932);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n7840, CK => CLK, Q => 
                           n15788, QN => n9937);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n7839, CK => CLK, Q => 
                           n15787, QN => n9942);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n7838, CK => CLK, Q => 
                           n15786, QN => n9947);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n7837, CK => CLK, Q => 
                           n15785, QN => n9952);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n7836, CK => CLK, Q => 
                           n15784, QN => n9957);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n7835, CK => CLK, Q => 
                           n15783, QN => n9962);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n7834, CK => CLK, Q => 
                           n15782, QN => n9967);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n7833, CK => CLK, Q => 
                           n15781, QN => n9972);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n7832, CK => CLK, Q => 
                           n15780, QN => n9977);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n7831, CK => CLK, Q => 
                           n15779, QN => n9982);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n7830, CK => CLK, Q => 
                           n15778, QN => n9987);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n7829, CK => CLK, Q => 
                           n15777, QN => n9992);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n7828, CK => CLK, Q => 
                           n15776, QN => n9997);
   REGISTERS_reg_1_63_inst : DFF_X1 port map( D => n7816, CK => CLK, Q => 
                           n15764, QN => n8969);
   REGISTERS_reg_1_62_inst : DFF_X1 port map( D => n7815, CK => CLK, Q => 
                           n15763, QN => n8974);
   REGISTERS_reg_1_61_inst : DFF_X1 port map( D => n7814, CK => CLK, Q => 
                           n15762, QN => n8979);
   REGISTERS_reg_1_60_inst : DFF_X1 port map( D => n7813, CK => CLK, Q => 
                           n15761, QN => n8984);
   REGISTERS_reg_1_59_inst : DFF_X1 port map( D => n7812, CK => CLK, Q => 
                           n15760, QN => n8989);
   REGISTERS_reg_1_58_inst : DFF_X1 port map( D => n7811, CK => CLK, Q => 
                           n15759, QN => n8994);
   REGISTERS_reg_1_57_inst : DFF_X1 port map( D => n7810, CK => CLK, Q => 
                           n15758, QN => n8999);
   REGISTERS_reg_1_56_inst : DFF_X1 port map( D => n7809, CK => CLK, Q => 
                           n15757, QN => n9004);
   REGISTERS_reg_1_55_inst : DFF_X1 port map( D => n7808, CK => CLK, Q => 
                           n15756, QN => n9009);
   REGISTERS_reg_1_54_inst : DFF_X1 port map( D => n7807, CK => CLK, Q => 
                           n15755, QN => n9014);
   REGISTERS_reg_1_53_inst : DFF_X1 port map( D => n7806, CK => CLK, Q => 
                           n15754, QN => n9019);
   REGISTERS_reg_1_52_inst : DFF_X1 port map( D => n7805, CK => CLK, Q => 
                           n15753, QN => n9024);
   REGISTERS_reg_1_51_inst : DFF_X1 port map( D => n7804, CK => CLK, Q => 
                           n15752, QN => n9029);
   REGISTERS_reg_1_50_inst : DFF_X1 port map( D => n7803, CK => CLK, Q => 
                           n15751, QN => n9034);
   REGISTERS_reg_1_49_inst : DFF_X1 port map( D => n7802, CK => CLK, Q => 
                           n15750, QN => n9039);
   REGISTERS_reg_1_48_inst : DFF_X1 port map( D => n7801, CK => CLK, Q => 
                           n15749, QN => n9044);
   REGISTERS_reg_1_47_inst : DFF_X1 port map( D => n7800, CK => CLK, Q => 
                           n15748, QN => n9049);
   REGISTERS_reg_1_46_inst : DFF_X1 port map( D => n7799, CK => CLK, Q => 
                           n15747, QN => n9054);
   REGISTERS_reg_1_45_inst : DFF_X1 port map( D => n7798, CK => CLK, Q => 
                           n15746, QN => n9059);
   REGISTERS_reg_1_44_inst : DFF_X1 port map( D => n7797, CK => CLK, Q => 
                           n15745, QN => n9064);
   REGISTERS_reg_1_43_inst : DFF_X1 port map( D => n7796, CK => CLK, Q => 
                           n15744, QN => n9069);
   REGISTERS_reg_1_42_inst : DFF_X1 port map( D => n7795, CK => CLK, Q => 
                           n15743, QN => n9074);
   REGISTERS_reg_1_41_inst : DFF_X1 port map( D => n7794, CK => CLK, Q => 
                           n15742, QN => n9079);
   REGISTERS_reg_1_40_inst : DFF_X1 port map( D => n7793, CK => CLK, Q => 
                           n15741, QN => n9084);
   REGISTERS_reg_1_39_inst : DFF_X1 port map( D => n7792, CK => CLK, Q => 
                           n15740, QN => n9089);
   REGISTERS_reg_1_38_inst : DFF_X1 port map( D => n7791, CK => CLK, Q => 
                           n15739, QN => n9094);
   REGISTERS_reg_1_37_inst : DFF_X1 port map( D => n7790, CK => CLK, Q => 
                           n15738, QN => n9099);
   REGISTERS_reg_1_36_inst : DFF_X1 port map( D => n7789, CK => CLK, Q => 
                           n15737, QN => n9104);
   REGISTERS_reg_1_35_inst : DFF_X1 port map( D => n7788, CK => CLK, Q => 
                           n15736, QN => n9109);
   REGISTERS_reg_1_34_inst : DFF_X1 port map( D => n7787, CK => CLK, Q => 
                           n15735, QN => n9114);
   REGISTERS_reg_1_33_inst : DFF_X1 port map( D => n7786, CK => CLK, Q => 
                           n15734, QN => n9119);
   REGISTERS_reg_1_32_inst : DFF_X1 port map( D => n7785, CK => CLK, Q => 
                           n15733, QN => n9124);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n7784, CK => CLK, Q => 
                           n15732, QN => n9129);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n7783, CK => CLK, Q => 
                           n15731, QN => n9134);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n7782, CK => CLK, Q => 
                           n15730, QN => n9139);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n7781, CK => CLK, Q => 
                           n15729, QN => n9144);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n7780, CK => CLK, Q => 
                           n15728, QN => n9149);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n7779, CK => CLK, Q => 
                           n15727, QN => n9154);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n7778, CK => CLK, Q => 
                           n15726, QN => n9159);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n7777, CK => CLK, Q => 
                           n15725, QN => n9164);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n7776, CK => CLK, Q => 
                           n15724, QN => n9169);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n7775, CK => CLK, Q => 
                           n15723, QN => n9174);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n7774, CK => CLK, Q => 
                           n15722, QN => n9179);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n7773, CK => CLK, Q => 
                           n15721, QN => n9184);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n7772, CK => CLK, Q => 
                           n15720, QN => n9189);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n7771, CK => CLK, Q => 
                           n15719, QN => n9194);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n7770, CK => CLK, Q => 
                           n15718, QN => n9199);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n7769, CK => CLK, Q => 
                           n15717, QN => n9204);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n7768, CK => CLK, Q => 
                           n15716, QN => n9209);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n7767, CK => CLK, Q => 
                           n15715, QN => n9214);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n7766, CK => CLK, Q => 
                           n15714, QN => n9219);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n7765, CK => CLK, Q => 
                           n15713, QN => n9224);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n7764, CK => CLK, Q => 
                           n15712, QN => n9229);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n7763, CK => CLK, Q => 
                           n15711, QN => n9234);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n7762, CK => CLK, Q => n15710
                           , QN => n9239);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n7761, CK => CLK, Q => n15709
                           , QN => n9244);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n7760, CK => CLK, Q => n15708
                           , QN => n9249);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n7759, CK => CLK, Q => n15707
                           , QN => n9254);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n7758, CK => CLK, Q => n15706
                           , QN => n9259);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n7757, CK => CLK, Q => n15705
                           , QN => n9264);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n7756, CK => CLK, Q => n15704
                           , QN => n9269);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n7755, CK => CLK, Q => n15703
                           , QN => n9274);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n7754, CK => CLK, Q => n15702
                           , QN => n9279);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n7753, CK => CLK, Q => n15701
                           , QN => n9284);
   REGISTERS_reg_4_63_inst : DFF_X1 port map( D => n7624, CK => CLK, Q => 
                           n15572, QN => n9738);
   REGISTERS_reg_4_62_inst : DFF_X1 port map( D => n7623, CK => CLK, Q => 
                           n15571, QN => n9743);
   REGISTERS_reg_4_61_inst : DFF_X1 port map( D => n7622, CK => CLK, Q => 
                           n15570, QN => n9748);
   REGISTERS_reg_4_60_inst : DFF_X1 port map( D => n7621, CK => CLK, Q => 
                           n15569, QN => n9753);
   REGISTERS_reg_4_59_inst : DFF_X1 port map( D => n7620, CK => CLK, Q => 
                           n15568, QN => n9758);
   REGISTERS_reg_4_58_inst : DFF_X1 port map( D => n7619, CK => CLK, Q => 
                           n15567, QN => n9763);
   REGISTERS_reg_4_57_inst : DFF_X1 port map( D => n7618, CK => CLK, Q => 
                           n15566, QN => n9768);
   REGISTERS_reg_4_56_inst : DFF_X1 port map( D => n7617, CK => CLK, Q => 
                           n15565, QN => n9773);
   REGISTERS_reg_4_55_inst : DFF_X1 port map( D => n7616, CK => CLK, Q => 
                           n15564, QN => n9778);
   REGISTERS_reg_4_54_inst : DFF_X1 port map( D => n7615, CK => CLK, Q => 
                           n15563, QN => n9783);
   REGISTERS_reg_4_53_inst : DFF_X1 port map( D => n7614, CK => CLK, Q => 
                           n15562, QN => n9788);
   REGISTERS_reg_4_52_inst : DFF_X1 port map( D => n7613, CK => CLK, Q => 
                           n15561, QN => n9793);
   REGISTERS_reg_4_51_inst : DFF_X1 port map( D => n7612, CK => CLK, Q => 
                           n15560, QN => n9798);
   REGISTERS_reg_4_50_inst : DFF_X1 port map( D => n7611, CK => CLK, Q => 
                           n15559, QN => n9803);
   REGISTERS_reg_4_49_inst : DFF_X1 port map( D => n7610, CK => CLK, Q => 
                           n15558, QN => n9808);
   REGISTERS_reg_4_48_inst : DFF_X1 port map( D => n7609, CK => CLK, Q => 
                           n15557, QN => n9813);
   REGISTERS_reg_4_47_inst : DFF_X1 port map( D => n7608, CK => CLK, Q => 
                           n15556, QN => n9818);
   REGISTERS_reg_4_46_inst : DFF_X1 port map( D => n7607, CK => CLK, Q => 
                           n15555, QN => n9823);
   REGISTERS_reg_4_45_inst : DFF_X1 port map( D => n7606, CK => CLK, Q => 
                           n15554, QN => n9828);
   REGISTERS_reg_4_44_inst : DFF_X1 port map( D => n7605, CK => CLK, Q => 
                           n15553, QN => n9833);
   REGISTERS_reg_4_43_inst : DFF_X1 port map( D => n7604, CK => CLK, Q => 
                           n15552, QN => n9838);
   REGISTERS_reg_4_42_inst : DFF_X1 port map( D => n7603, CK => CLK, Q => 
                           n15551, QN => n9843);
   REGISTERS_reg_4_41_inst : DFF_X1 port map( D => n7602, CK => CLK, Q => 
                           n15550, QN => n9848);
   REGISTERS_reg_4_40_inst : DFF_X1 port map( D => n7601, CK => CLK, Q => 
                           n15549, QN => n9853);
   REGISTERS_reg_4_39_inst : DFF_X1 port map( D => n7600, CK => CLK, Q => 
                           n15548, QN => n9858);
   REGISTERS_reg_4_38_inst : DFF_X1 port map( D => n7599, CK => CLK, Q => 
                           n15547, QN => n9863);
   REGISTERS_reg_4_37_inst : DFF_X1 port map( D => n7598, CK => CLK, Q => 
                           n15546, QN => n9868);
   REGISTERS_reg_4_36_inst : DFF_X1 port map( D => n7597, CK => CLK, Q => 
                           n15545, QN => n9873);
   REGISTERS_reg_4_35_inst : DFF_X1 port map( D => n7596, CK => CLK, Q => 
                           n15544, QN => n9878);
   REGISTERS_reg_4_34_inst : DFF_X1 port map( D => n7595, CK => CLK, Q => 
                           n15543, QN => n9883);
   REGISTERS_reg_4_33_inst : DFF_X1 port map( D => n7594, CK => CLK, Q => 
                           n15542, QN => n9888);
   REGISTERS_reg_4_32_inst : DFF_X1 port map( D => n7593, CK => CLK, Q => 
                           n15541, QN => n9893);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n7592, CK => CLK, Q => 
                           n15540, QN => n9898);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n7591, CK => CLK, Q => 
                           n15539, QN => n9903);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n7590, CK => CLK, Q => 
                           n15538, QN => n9908);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n7589, CK => CLK, Q => 
                           n15537, QN => n9913);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n7588, CK => CLK, Q => 
                           n15536, QN => n9918);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n7587, CK => CLK, Q => 
                           n15535, QN => n9923);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n7586, CK => CLK, Q => 
                           n15534, QN => n9928);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n7585, CK => CLK, Q => 
                           n15533, QN => n9933);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n7584, CK => CLK, Q => 
                           n15532, QN => n9938);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n7583, CK => CLK, Q => 
                           n15531, QN => n9943);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n7582, CK => CLK, Q => 
                           n15530, QN => n9948);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n7581, CK => CLK, Q => 
                           n15529, QN => n9953);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n7580, CK => CLK, Q => 
                           n15528, QN => n9958);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n7579, CK => CLK, Q => 
                           n15527, QN => n9963);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n7578, CK => CLK, Q => 
                           n15526, QN => n9968);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n7577, CK => CLK, Q => 
                           n15525, QN => n9973);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n7576, CK => CLK, Q => 
                           n15524, QN => n9978);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n7575, CK => CLK, Q => 
                           n15523, QN => n9983);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n7574, CK => CLK, Q => 
                           n15522, QN => n9988);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n7573, CK => CLK, Q => 
                           n15521, QN => n9993);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n7572, CK => CLK, Q => 
                           n15520, QN => n9998);
   REGISTERS_reg_5_63_inst : DFF_X1 port map( D => n7560, CK => CLK, Q => 
                           n15508, QN => n8970);
   REGISTERS_reg_5_62_inst : DFF_X1 port map( D => n7559, CK => CLK, Q => 
                           n15507, QN => n8975);
   REGISTERS_reg_5_61_inst : DFF_X1 port map( D => n7558, CK => CLK, Q => 
                           n15506, QN => n8980);
   REGISTERS_reg_5_60_inst : DFF_X1 port map( D => n7557, CK => CLK, Q => 
                           n15505, QN => n8985);
   REGISTERS_reg_5_59_inst : DFF_X1 port map( D => n7556, CK => CLK, Q => 
                           n15504, QN => n8990);
   REGISTERS_reg_5_58_inst : DFF_X1 port map( D => n7555, CK => CLK, Q => 
                           n15503, QN => n8995);
   REGISTERS_reg_5_57_inst : DFF_X1 port map( D => n7554, CK => CLK, Q => 
                           n15502, QN => n9000);
   REGISTERS_reg_5_56_inst : DFF_X1 port map( D => n7553, CK => CLK, Q => 
                           n15501, QN => n9005);
   REGISTERS_reg_5_55_inst : DFF_X1 port map( D => n7552, CK => CLK, Q => 
                           n15500, QN => n9010);
   REGISTERS_reg_5_54_inst : DFF_X1 port map( D => n7551, CK => CLK, Q => 
                           n15499, QN => n9015);
   REGISTERS_reg_5_53_inst : DFF_X1 port map( D => n7550, CK => CLK, Q => 
                           n15498, QN => n9020);
   REGISTERS_reg_5_52_inst : DFF_X1 port map( D => n7549, CK => CLK, Q => 
                           n15497, QN => n9025);
   REGISTERS_reg_5_51_inst : DFF_X1 port map( D => n7548, CK => CLK, Q => 
                           n15496, QN => n9030);
   REGISTERS_reg_5_50_inst : DFF_X1 port map( D => n7547, CK => CLK, Q => 
                           n15495, QN => n9035);
   REGISTERS_reg_5_49_inst : DFF_X1 port map( D => n7546, CK => CLK, Q => 
                           n15494, QN => n9040);
   REGISTERS_reg_5_48_inst : DFF_X1 port map( D => n7545, CK => CLK, Q => 
                           n15493, QN => n9045);
   REGISTERS_reg_5_47_inst : DFF_X1 port map( D => n7544, CK => CLK, Q => 
                           n15492, QN => n9050);
   REGISTERS_reg_5_46_inst : DFF_X1 port map( D => n7543, CK => CLK, Q => 
                           n15491, QN => n9055);
   REGISTERS_reg_5_45_inst : DFF_X1 port map( D => n7542, CK => CLK, Q => 
                           n15490, QN => n9060);
   REGISTERS_reg_5_44_inst : DFF_X1 port map( D => n7541, CK => CLK, Q => 
                           n15489, QN => n9065);
   REGISTERS_reg_5_43_inst : DFF_X1 port map( D => n7540, CK => CLK, Q => 
                           n15488, QN => n9070);
   REGISTERS_reg_5_42_inst : DFF_X1 port map( D => n7539, CK => CLK, Q => 
                           n15487, QN => n9075);
   REGISTERS_reg_5_41_inst : DFF_X1 port map( D => n7538, CK => CLK, Q => 
                           n15486, QN => n9080);
   REGISTERS_reg_5_40_inst : DFF_X1 port map( D => n7537, CK => CLK, Q => 
                           n15485, QN => n9085);
   REGISTERS_reg_5_39_inst : DFF_X1 port map( D => n7536, CK => CLK, Q => 
                           n15484, QN => n9090);
   REGISTERS_reg_5_38_inst : DFF_X1 port map( D => n7535, CK => CLK, Q => 
                           n15483, QN => n9095);
   REGISTERS_reg_5_37_inst : DFF_X1 port map( D => n7534, CK => CLK, Q => 
                           n15482, QN => n9100);
   REGISTERS_reg_5_36_inst : DFF_X1 port map( D => n7533, CK => CLK, Q => 
                           n15481, QN => n9105);
   REGISTERS_reg_5_35_inst : DFF_X1 port map( D => n7532, CK => CLK, Q => 
                           n15480, QN => n9110);
   REGISTERS_reg_5_34_inst : DFF_X1 port map( D => n7531, CK => CLK, Q => 
                           n15479, QN => n9115);
   REGISTERS_reg_5_33_inst : DFF_X1 port map( D => n7530, CK => CLK, Q => 
                           n15478, QN => n9120);
   REGISTERS_reg_5_32_inst : DFF_X1 port map( D => n7529, CK => CLK, Q => 
                           n15477, QN => n9125);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n7528, CK => CLK, Q => 
                           n15476, QN => n9130);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n7527, CK => CLK, Q => 
                           n15475, QN => n9135);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n7526, CK => CLK, Q => 
                           n15474, QN => n9140);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n7525, CK => CLK, Q => 
                           n15473, QN => n9145);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n7524, CK => CLK, Q => 
                           n15472, QN => n9150);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n7523, CK => CLK, Q => 
                           n15471, QN => n9155);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n7522, CK => CLK, Q => 
                           n15470, QN => n9160);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n7521, CK => CLK, Q => 
                           n15469, QN => n9165);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n7520, CK => CLK, Q => 
                           n15468, QN => n9170);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n7519, CK => CLK, Q => 
                           n15467, QN => n9175);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n7518, CK => CLK, Q => 
                           n15466, QN => n9180);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n7517, CK => CLK, Q => 
                           n15465, QN => n9185);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n7516, CK => CLK, Q => 
                           n15464, QN => n9190);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n7515, CK => CLK, Q => 
                           n15463, QN => n9195);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n7514, CK => CLK, Q => 
                           n15462, QN => n9200);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n7513, CK => CLK, Q => 
                           n15461, QN => n9205);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n7512, CK => CLK, Q => 
                           n15460, QN => n9210);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n7511, CK => CLK, Q => 
                           n15459, QN => n9215);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n7510, CK => CLK, Q => 
                           n15458, QN => n9220);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n7509, CK => CLK, Q => 
                           n15457, QN => n9225);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n7508, CK => CLK, Q => 
                           n15456, QN => n9230);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n7507, CK => CLK, Q => 
                           n15455, QN => n9235);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n7506, CK => CLK, Q => n15454
                           , QN => n9240);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n7505, CK => CLK, Q => n15453
                           , QN => n9245);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n7504, CK => CLK, Q => n15452
                           , QN => n9250);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n7503, CK => CLK, Q => n15451
                           , QN => n9255);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n7502, CK => CLK, Q => n15450
                           , QN => n9260);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n7501, CK => CLK, Q => n15449
                           , QN => n9265);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n7500, CK => CLK, Q => n15448
                           , QN => n9270);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n7499, CK => CLK, Q => n15447
                           , QN => n9275);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n7498, CK => CLK, Q => n15446
                           , QN => n9280);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n7497, CK => CLK, Q => n15445
                           , QN => n9285);
   REGISTERS_reg_10_63_inst : DFF_X1 port map( D => n7240, CK => CLK, Q => 
                           n15188, QN => n9739);
   REGISTERS_reg_10_62_inst : DFF_X1 port map( D => n7239, CK => CLK, Q => 
                           n15187, QN => n9744);
   REGISTERS_reg_10_61_inst : DFF_X1 port map( D => n7238, CK => CLK, Q => 
                           n15186, QN => n9749);
   REGISTERS_reg_10_60_inst : DFF_X1 port map( D => n7237, CK => CLK, Q => 
                           n15185, QN => n9754);
   REGISTERS_reg_10_59_inst : DFF_X1 port map( D => n7236, CK => CLK, Q => 
                           n15184, QN => n9759);
   REGISTERS_reg_10_58_inst : DFF_X1 port map( D => n7235, CK => CLK, Q => 
                           n15183, QN => n9764);
   REGISTERS_reg_10_57_inst : DFF_X1 port map( D => n7234, CK => CLK, Q => 
                           n15182, QN => n9769);
   REGISTERS_reg_10_56_inst : DFF_X1 port map( D => n7233, CK => CLK, Q => 
                           n15181, QN => n9774);
   REGISTERS_reg_10_55_inst : DFF_X1 port map( D => n7232, CK => CLK, Q => 
                           n15180, QN => n9779);
   REGISTERS_reg_10_54_inst : DFF_X1 port map( D => n7231, CK => CLK, Q => 
                           n15179, QN => n9784);
   REGISTERS_reg_10_53_inst : DFF_X1 port map( D => n7230, CK => CLK, Q => 
                           n15178, QN => n9789);
   REGISTERS_reg_10_52_inst : DFF_X1 port map( D => n7229, CK => CLK, Q => 
                           n15177, QN => n9794);
   REGISTERS_reg_10_51_inst : DFF_X1 port map( D => n7228, CK => CLK, Q => 
                           n15176, QN => n9799);
   REGISTERS_reg_10_50_inst : DFF_X1 port map( D => n7227, CK => CLK, Q => 
                           n15175, QN => n9804);
   REGISTERS_reg_10_49_inst : DFF_X1 port map( D => n7226, CK => CLK, Q => 
                           n15174, QN => n9809);
   REGISTERS_reg_10_48_inst : DFF_X1 port map( D => n7225, CK => CLK, Q => 
                           n15173, QN => n9814);
   REGISTERS_reg_10_47_inst : DFF_X1 port map( D => n7224, CK => CLK, Q => 
                           n15172, QN => n9819);
   REGISTERS_reg_10_46_inst : DFF_X1 port map( D => n7223, CK => CLK, Q => 
                           n15171, QN => n9824);
   REGISTERS_reg_10_45_inst : DFF_X1 port map( D => n7222, CK => CLK, Q => 
                           n15170, QN => n9829);
   REGISTERS_reg_10_44_inst : DFF_X1 port map( D => n7221, CK => CLK, Q => 
                           n15169, QN => n9834);
   REGISTERS_reg_10_43_inst : DFF_X1 port map( D => n7220, CK => CLK, Q => 
                           n15168, QN => n9839);
   REGISTERS_reg_10_42_inst : DFF_X1 port map( D => n7219, CK => CLK, Q => 
                           n15167, QN => n9844);
   REGISTERS_reg_10_41_inst : DFF_X1 port map( D => n7218, CK => CLK, Q => 
                           n15166, QN => n9849);
   REGISTERS_reg_10_40_inst : DFF_X1 port map( D => n7217, CK => CLK, Q => 
                           n15165, QN => n9854);
   REGISTERS_reg_10_39_inst : DFF_X1 port map( D => n7216, CK => CLK, Q => 
                           n15164, QN => n9859);
   REGISTERS_reg_10_38_inst : DFF_X1 port map( D => n7215, CK => CLK, Q => 
                           n15163, QN => n9864);
   REGISTERS_reg_10_37_inst : DFF_X1 port map( D => n7214, CK => CLK, Q => 
                           n15162, QN => n9869);
   REGISTERS_reg_10_36_inst : DFF_X1 port map( D => n7213, CK => CLK, Q => 
                           n15161, QN => n9874);
   REGISTERS_reg_10_35_inst : DFF_X1 port map( D => n7212, CK => CLK, Q => 
                           n15160, QN => n9879);
   REGISTERS_reg_10_34_inst : DFF_X1 port map( D => n7211, CK => CLK, Q => 
                           n15159, QN => n9884);
   REGISTERS_reg_10_33_inst : DFF_X1 port map( D => n7210, CK => CLK, Q => 
                           n15158, QN => n9889);
   REGISTERS_reg_10_32_inst : DFF_X1 port map( D => n7209, CK => CLK, Q => 
                           n15157, QN => n9894);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n7208, CK => CLK, Q => 
                           n15156, QN => n9899);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n7207, CK => CLK, Q => 
                           n15155, QN => n9904);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n7206, CK => CLK, Q => 
                           n15154, QN => n9909);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n7205, CK => CLK, Q => 
                           n15153, QN => n9914);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n7204, CK => CLK, Q => 
                           n15152, QN => n9919);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n7203, CK => CLK, Q => 
                           n15151, QN => n9924);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n7202, CK => CLK, Q => 
                           n15150, QN => n9929);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n7201, CK => CLK, Q => 
                           n15149, QN => n9934);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n7200, CK => CLK, Q => 
                           n15148, QN => n9939);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n7199, CK => CLK, Q => 
                           n15147, QN => n9944);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n7198, CK => CLK, Q => 
                           n15146, QN => n9949);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n7197, CK => CLK, Q => 
                           n15145, QN => n9954);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n7196, CK => CLK, Q => 
                           n15144, QN => n9959);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n7195, CK => CLK, Q => 
                           n15143, QN => n9964);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n7194, CK => CLK, Q => 
                           n15142, QN => n9969);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n7193, CK => CLK, Q => 
                           n15141, QN => n9974);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n7192, CK => CLK, Q => 
                           n15140, QN => n9979);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n7191, CK => CLK, Q => 
                           n15139, QN => n9984);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n7190, CK => CLK, Q => 
                           n15138, QN => n9989);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n7189, CK => CLK, Q => 
                           n15137, QN => n9994);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n7188, CK => CLK, Q => 
                           n15136, QN => n9999);
   REGISTERS_reg_11_63_inst : DFF_X1 port map( D => n7176, CK => CLK, Q => 
                           n15124, QN => n8971);
   REGISTERS_reg_11_62_inst : DFF_X1 port map( D => n7175, CK => CLK, Q => 
                           n15123, QN => n8976);
   REGISTERS_reg_11_61_inst : DFF_X1 port map( D => n7174, CK => CLK, Q => 
                           n15122, QN => n8981);
   REGISTERS_reg_11_60_inst : DFF_X1 port map( D => n7173, CK => CLK, Q => 
                           n15121, QN => n8986);
   REGISTERS_reg_11_59_inst : DFF_X1 port map( D => n7172, CK => CLK, Q => 
                           n15120, QN => n8991);
   REGISTERS_reg_11_58_inst : DFF_X1 port map( D => n7171, CK => CLK, Q => 
                           n15119, QN => n8996);
   REGISTERS_reg_11_57_inst : DFF_X1 port map( D => n7170, CK => CLK, Q => 
                           n15118, QN => n9001);
   REGISTERS_reg_11_56_inst : DFF_X1 port map( D => n7169, CK => CLK, Q => 
                           n15117, QN => n9006);
   REGISTERS_reg_11_55_inst : DFF_X1 port map( D => n7168, CK => CLK, Q => 
                           n15116, QN => n9011);
   REGISTERS_reg_11_54_inst : DFF_X1 port map( D => n7167, CK => CLK, Q => 
                           n15115, QN => n9016);
   REGISTERS_reg_11_53_inst : DFF_X1 port map( D => n7166, CK => CLK, Q => 
                           n15114, QN => n9021);
   REGISTERS_reg_11_52_inst : DFF_X1 port map( D => n7165, CK => CLK, Q => 
                           n15113, QN => n9026);
   REGISTERS_reg_11_51_inst : DFF_X1 port map( D => n7164, CK => CLK, Q => 
                           n15112, QN => n9031);
   REGISTERS_reg_11_50_inst : DFF_X1 port map( D => n7163, CK => CLK, Q => 
                           n15111, QN => n9036);
   REGISTERS_reg_11_49_inst : DFF_X1 port map( D => n7162, CK => CLK, Q => 
                           n15110, QN => n9041);
   REGISTERS_reg_11_48_inst : DFF_X1 port map( D => n7161, CK => CLK, Q => 
                           n15109, QN => n9046);
   REGISTERS_reg_11_47_inst : DFF_X1 port map( D => n7160, CK => CLK, Q => 
                           n15108, QN => n9051);
   REGISTERS_reg_11_46_inst : DFF_X1 port map( D => n7159, CK => CLK, Q => 
                           n15107, QN => n9056);
   REGISTERS_reg_11_45_inst : DFF_X1 port map( D => n7158, CK => CLK, Q => 
                           n15106, QN => n9061);
   REGISTERS_reg_11_44_inst : DFF_X1 port map( D => n7157, CK => CLK, Q => 
                           n15105, QN => n9066);
   REGISTERS_reg_11_43_inst : DFF_X1 port map( D => n7156, CK => CLK, Q => 
                           n15104, QN => n9071);
   REGISTERS_reg_11_42_inst : DFF_X1 port map( D => n7155, CK => CLK, Q => 
                           n15103, QN => n9076);
   REGISTERS_reg_11_41_inst : DFF_X1 port map( D => n7154, CK => CLK, Q => 
                           n15102, QN => n9081);
   REGISTERS_reg_11_40_inst : DFF_X1 port map( D => n7153, CK => CLK, Q => 
                           n15101, QN => n9086);
   REGISTERS_reg_11_39_inst : DFF_X1 port map( D => n7152, CK => CLK, Q => 
                           n15100, QN => n9091);
   REGISTERS_reg_11_38_inst : DFF_X1 port map( D => n7151, CK => CLK, Q => 
                           n15099, QN => n9096);
   REGISTERS_reg_11_37_inst : DFF_X1 port map( D => n7150, CK => CLK, Q => 
                           n15098, QN => n9101);
   REGISTERS_reg_11_36_inst : DFF_X1 port map( D => n7149, CK => CLK, Q => 
                           n15097, QN => n9106);
   REGISTERS_reg_11_35_inst : DFF_X1 port map( D => n7148, CK => CLK, Q => 
                           n15096, QN => n9111);
   REGISTERS_reg_11_34_inst : DFF_X1 port map( D => n7147, CK => CLK, Q => 
                           n15095, QN => n9116);
   REGISTERS_reg_11_33_inst : DFF_X1 port map( D => n7146, CK => CLK, Q => 
                           n15094, QN => n9121);
   REGISTERS_reg_11_32_inst : DFF_X1 port map( D => n7145, CK => CLK, Q => 
                           n15093, QN => n9126);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n7144, CK => CLK, Q => 
                           n15092, QN => n9131);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n7143, CK => CLK, Q => 
                           n15091, QN => n9136);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n7142, CK => CLK, Q => 
                           n15090, QN => n9141);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n7141, CK => CLK, Q => 
                           n15089, QN => n9146);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n7140, CK => CLK, Q => 
                           n15088, QN => n9151);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n7139, CK => CLK, Q => 
                           n15087, QN => n9156);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n7138, CK => CLK, Q => 
                           n15086, QN => n9161);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n7137, CK => CLK, Q => 
                           n15085, QN => n9166);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n7136, CK => CLK, Q => 
                           n15084, QN => n9171);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n7135, CK => CLK, Q => 
                           n15083, QN => n9176);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n7134, CK => CLK, Q => 
                           n15082, QN => n9181);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n7133, CK => CLK, Q => 
                           n15081, QN => n9186);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n7132, CK => CLK, Q => 
                           n15080, QN => n9191);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n7131, CK => CLK, Q => 
                           n15079, QN => n9196);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n7130, CK => CLK, Q => 
                           n15078, QN => n9201);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n7129, CK => CLK, Q => 
                           n15077, QN => n9206);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n7128, CK => CLK, Q => 
                           n15076, QN => n9211);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n7127, CK => CLK, Q => 
                           n15075, QN => n9216);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n7126, CK => CLK, Q => 
                           n15074, QN => n9221);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n7125, CK => CLK, Q => 
                           n15073, QN => n9226);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n7124, CK => CLK, Q => 
                           n15072, QN => n9231);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n7123, CK => CLK, Q => 
                           n15071, QN => n9236);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n7122, CK => CLK, Q => 
                           n15070, QN => n9241);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n7121, CK => CLK, Q => 
                           n15069, QN => n9246);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n7120, CK => CLK, Q => 
                           n15068, QN => n9251);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n7119, CK => CLK, Q => 
                           n15067, QN => n9256);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n7118, CK => CLK, Q => 
                           n15066, QN => n9261);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n7117, CK => CLK, Q => 
                           n15065, QN => n9266);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n7116, CK => CLK, Q => 
                           n15064, QN => n9271);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n7115, CK => CLK, Q => 
                           n15063, QN => n9276);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n7114, CK => CLK, Q => 
                           n15062, QN => n9281);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n7113, CK => CLK, Q => 
                           n15061, QN => n9286);
   REGISTERS_reg_15_63_inst : DFF_X1 port map( D => n6920, CK => CLK, Q => 
                           n29827, QN => n9609);
   REGISTERS_reg_15_62_inst : DFF_X1 port map( D => n6919, CK => CLK, Q => 
                           n29826, QN => n9610);
   REGISTERS_reg_15_61_inst : DFF_X1 port map( D => n6918, CK => CLK, Q => 
                           n29825, QN => n9611);
   REGISTERS_reg_15_60_inst : DFF_X1 port map( D => n6917, CK => CLK, Q => 
                           n29824, QN => n9612);
   REGISTERS_reg_15_59_inst : DFF_X1 port map( D => n6916, CK => CLK, Q => 
                           n29823, QN => n9613);
   REGISTERS_reg_15_58_inst : DFF_X1 port map( D => n6915, CK => CLK, Q => 
                           n29822, QN => n9614);
   REGISTERS_reg_15_57_inst : DFF_X1 port map( D => n6914, CK => CLK, Q => 
                           n29821, QN => n9615);
   REGISTERS_reg_15_56_inst : DFF_X1 port map( D => n6913, CK => CLK, Q => 
                           n29820, QN => n9616);
   REGISTERS_reg_15_55_inst : DFF_X1 port map( D => n6912, CK => CLK, Q => 
                           n29819, QN => n9617);
   REGISTERS_reg_15_54_inst : DFF_X1 port map( D => n6911, CK => CLK, Q => 
                           n29818, QN => n9618);
   REGISTERS_reg_15_53_inst : DFF_X1 port map( D => n6910, CK => CLK, Q => 
                           n29817, QN => n9619);
   REGISTERS_reg_15_52_inst : DFF_X1 port map( D => n6909, CK => CLK, Q => 
                           n29816, QN => n9620);
   REGISTERS_reg_15_51_inst : DFF_X1 port map( D => n6908, CK => CLK, Q => 
                           n29815, QN => n9621);
   REGISTERS_reg_15_50_inst : DFF_X1 port map( D => n6907, CK => CLK, Q => 
                           n29814, QN => n9622);
   REGISTERS_reg_15_49_inst : DFF_X1 port map( D => n6906, CK => CLK, Q => 
                           n29813, QN => n9623);
   REGISTERS_reg_15_48_inst : DFF_X1 port map( D => n6905, CK => CLK, Q => 
                           n29812, QN => n9624);
   REGISTERS_reg_15_47_inst : DFF_X1 port map( D => n6904, CK => CLK, Q => 
                           n29811, QN => n9625);
   REGISTERS_reg_15_46_inst : DFF_X1 port map( D => n6903, CK => CLK, Q => 
                           n29810, QN => n9626);
   REGISTERS_reg_15_45_inst : DFF_X1 port map( D => n6902, CK => CLK, Q => 
                           n29809, QN => n9627);
   REGISTERS_reg_15_44_inst : DFF_X1 port map( D => n6901, CK => CLK, Q => 
                           n29808, QN => n9628);
   REGISTERS_reg_15_43_inst : DFF_X1 port map( D => n6900, CK => CLK, Q => 
                           n29807, QN => n9629);
   REGISTERS_reg_15_42_inst : DFF_X1 port map( D => n6899, CK => CLK, Q => 
                           n29806, QN => n9630);
   REGISTERS_reg_15_41_inst : DFF_X1 port map( D => n6898, CK => CLK, Q => 
                           n29805, QN => n9631);
   REGISTERS_reg_15_40_inst : DFF_X1 port map( D => n6897, CK => CLK, Q => 
                           n29804, QN => n9632);
   REGISTERS_reg_15_39_inst : DFF_X1 port map( D => n6896, CK => CLK, Q => 
                           n29803, QN => n9633);
   REGISTERS_reg_15_38_inst : DFF_X1 port map( D => n6895, CK => CLK, Q => 
                           n29802, QN => n9634);
   REGISTERS_reg_15_37_inst : DFF_X1 port map( D => n6894, CK => CLK, Q => 
                           n29801, QN => n9635);
   REGISTERS_reg_15_36_inst : DFF_X1 port map( D => n6893, CK => CLK, Q => 
                           n29800, QN => n9636);
   REGISTERS_reg_15_35_inst : DFF_X1 port map( D => n6892, CK => CLK, Q => 
                           n29799, QN => n9637);
   REGISTERS_reg_15_34_inst : DFF_X1 port map( D => n6891, CK => CLK, Q => 
                           n29798, QN => n9638);
   REGISTERS_reg_15_33_inst : DFF_X1 port map( D => n6890, CK => CLK, Q => 
                           n29797, QN => n9639);
   REGISTERS_reg_15_32_inst : DFF_X1 port map( D => n6889, CK => CLK, Q => 
                           n29796, QN => n9640);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n6888, CK => CLK, Q => 
                           n29795, QN => n9641);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n6887, CK => CLK, Q => 
                           n29794, QN => n9642);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n6886, CK => CLK, Q => 
                           n29793, QN => n9643);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n6885, CK => CLK, Q => 
                           n29792, QN => n9644);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n6884, CK => CLK, Q => 
                           n29791, QN => n9645);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n6883, CK => CLK, Q => 
                           n29790, QN => n9646);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n6882, CK => CLK, Q => 
                           n29789, QN => n9647);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n6881, CK => CLK, Q => 
                           n29788, QN => n9648);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n6880, CK => CLK, Q => 
                           n29787, QN => n9649);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n6879, CK => CLK, Q => 
                           n29786, QN => n9650);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n6878, CK => CLK, Q => 
                           n29785, QN => n9651);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n6877, CK => CLK, Q => 
                           n29784, QN => n9652);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n6876, CK => CLK, Q => 
                           n29783, QN => n9653);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n6875, CK => CLK, Q => 
                           n29782, QN => n9654);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n6874, CK => CLK, Q => 
                           n29781, QN => n9655);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n6873, CK => CLK, Q => 
                           n29780, QN => n9656);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n6872, CK => CLK, Q => 
                           n29779, QN => n9657);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n6871, CK => CLK, Q => 
                           n29778, QN => n9658);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n6870, CK => CLK, Q => 
                           n29777, QN => n9659);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n6869, CK => CLK, Q => 
                           n29776, QN => n9660);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n6868, CK => CLK, Q => 
                           n29775, QN => n9661);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n6867, CK => CLK, Q => 
                           n29774, QN => n9662);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n6866, CK => CLK, Q => 
                           n29773, QN => n9663);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n6865, CK => CLK, Q => 
                           n29772, QN => n9664);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n6864, CK => CLK, Q => 
                           n29771, QN => n9665);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n6863, CK => CLK, Q => 
                           n29770, QN => n9666);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n6862, CK => CLK, Q => 
                           n29769, QN => n9667);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n6861, CK => CLK, Q => 
                           n29768, QN => n9668);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n6860, CK => CLK, Q => 
                           n29767, QN => n9669);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n6859, CK => CLK, Q => 
                           n29766, QN => n9670);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n6858, CK => CLK, Q => 
                           n29765, QN => n9671);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n6857, CK => CLK, Q => 
                           n29764, QN => n9672);
   REGISTERS_reg_18_63_inst : DFF_X1 port map( D => n6728, CK => CLK, Q => 
                           n14676, QN => n9741);
   REGISTERS_reg_18_62_inst : DFF_X1 port map( D => n6727, CK => CLK, Q => 
                           n14675, QN => n9746);
   REGISTERS_reg_18_61_inst : DFF_X1 port map( D => n6726, CK => CLK, Q => 
                           n14674, QN => n9751);
   REGISTERS_reg_18_60_inst : DFF_X1 port map( D => n6725, CK => CLK, Q => 
                           n14673, QN => n9756);
   REGISTERS_reg_18_59_inst : DFF_X1 port map( D => n6724, CK => CLK, Q => 
                           n14672, QN => n9761);
   REGISTERS_reg_18_58_inst : DFF_X1 port map( D => n6723, CK => CLK, Q => 
                           n14671, QN => n9766);
   REGISTERS_reg_18_57_inst : DFF_X1 port map( D => n6722, CK => CLK, Q => 
                           n14670, QN => n9771);
   REGISTERS_reg_18_56_inst : DFF_X1 port map( D => n6721, CK => CLK, Q => 
                           n14669, QN => n9776);
   REGISTERS_reg_18_55_inst : DFF_X1 port map( D => n6720, CK => CLK, Q => 
                           n14668, QN => n9781);
   REGISTERS_reg_18_54_inst : DFF_X1 port map( D => n6719, CK => CLK, Q => 
                           n14667, QN => n9786);
   REGISTERS_reg_18_53_inst : DFF_X1 port map( D => n6718, CK => CLK, Q => 
                           n14666, QN => n9791);
   REGISTERS_reg_18_52_inst : DFF_X1 port map( D => n6717, CK => CLK, Q => 
                           n14665, QN => n9796);
   REGISTERS_reg_18_51_inst : DFF_X1 port map( D => n6716, CK => CLK, Q => 
                           n14664, QN => n9801);
   REGISTERS_reg_18_50_inst : DFF_X1 port map( D => n6715, CK => CLK, Q => 
                           n14663, QN => n9806);
   REGISTERS_reg_18_49_inst : DFF_X1 port map( D => n6714, CK => CLK, Q => 
                           n14662, QN => n9811);
   REGISTERS_reg_18_48_inst : DFF_X1 port map( D => n6713, CK => CLK, Q => 
                           n14661, QN => n9816);
   REGISTERS_reg_18_47_inst : DFF_X1 port map( D => n6712, CK => CLK, Q => 
                           n14660, QN => n9821);
   REGISTERS_reg_18_46_inst : DFF_X1 port map( D => n6711, CK => CLK, Q => 
                           n14659, QN => n9826);
   REGISTERS_reg_18_45_inst : DFF_X1 port map( D => n6710, CK => CLK, Q => 
                           n14658, QN => n9831);
   REGISTERS_reg_18_44_inst : DFF_X1 port map( D => n6709, CK => CLK, Q => 
                           n14657, QN => n9836);
   REGISTERS_reg_18_43_inst : DFF_X1 port map( D => n6708, CK => CLK, Q => 
                           n14656, QN => n9841);
   REGISTERS_reg_18_42_inst : DFF_X1 port map( D => n6707, CK => CLK, Q => 
                           n14655, QN => n9846);
   REGISTERS_reg_18_41_inst : DFF_X1 port map( D => n6706, CK => CLK, Q => 
                           n14654, QN => n9851);
   REGISTERS_reg_18_40_inst : DFF_X1 port map( D => n6705, CK => CLK, Q => 
                           n14653, QN => n9856);
   REGISTERS_reg_18_39_inst : DFF_X1 port map( D => n6704, CK => CLK, Q => 
                           n14652, QN => n9861);
   REGISTERS_reg_18_38_inst : DFF_X1 port map( D => n6703, CK => CLK, Q => 
                           n14651, QN => n9866);
   REGISTERS_reg_18_37_inst : DFF_X1 port map( D => n6702, CK => CLK, Q => 
                           n14650, QN => n9871);
   REGISTERS_reg_18_36_inst : DFF_X1 port map( D => n6701, CK => CLK, Q => 
                           n14649, QN => n9876);
   REGISTERS_reg_18_35_inst : DFF_X1 port map( D => n6700, CK => CLK, Q => 
                           n14648, QN => n9881);
   REGISTERS_reg_18_34_inst : DFF_X1 port map( D => n6699, CK => CLK, Q => 
                           n14647, QN => n9886);
   REGISTERS_reg_18_33_inst : DFF_X1 port map( D => n6698, CK => CLK, Q => 
                           n14646, QN => n9891);
   REGISTERS_reg_18_32_inst : DFF_X1 port map( D => n6697, CK => CLK, Q => 
                           n14645, QN => n9896);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n6696, CK => CLK, Q => 
                           n14644, QN => n9901);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n6695, CK => CLK, Q => 
                           n14643, QN => n9906);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n6694, CK => CLK, Q => 
                           n14642, QN => n9911);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n6693, CK => CLK, Q => 
                           n14641, QN => n9916);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n6692, CK => CLK, Q => 
                           n14640, QN => n9921);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n6691, CK => CLK, Q => 
                           n14639, QN => n9926);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n6690, CK => CLK, Q => 
                           n14638, QN => n9931);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n6689, CK => CLK, Q => 
                           n14637, QN => n9936);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n6688, CK => CLK, Q => 
                           n14636, QN => n9941);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n6687, CK => CLK, Q => 
                           n14635, QN => n9946);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n6686, CK => CLK, Q => 
                           n14634, QN => n9951);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n6685, CK => CLK, Q => 
                           n14633, QN => n9956);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n6684, CK => CLK, Q => 
                           n14632, QN => n9961);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n6683, CK => CLK, Q => 
                           n14631, QN => n9966);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n6682, CK => CLK, Q => 
                           n14630, QN => n9971);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n6681, CK => CLK, Q => 
                           n14629, QN => n9976);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n6680, CK => CLK, Q => 
                           n14628, QN => n9981);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n6679, CK => CLK, Q => 
                           n14627, QN => n9986);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n6678, CK => CLK, Q => 
                           n14626, QN => n9991);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n6677, CK => CLK, Q => 
                           n14625, QN => n9996);
   REGISTERS_reg_19_63_inst : DFF_X1 port map( D => n6664, CK => CLK, Q => 
                           n14612, QN => n8973);
   REGISTERS_reg_19_62_inst : DFF_X1 port map( D => n6663, CK => CLK, Q => 
                           n14611, QN => n8978);
   REGISTERS_reg_19_61_inst : DFF_X1 port map( D => n6662, CK => CLK, Q => 
                           n14610, QN => n8983);
   REGISTERS_reg_19_60_inst : DFF_X1 port map( D => n6661, CK => CLK, Q => 
                           n14609, QN => n8988);
   REGISTERS_reg_19_59_inst : DFF_X1 port map( D => n6660, CK => CLK, Q => 
                           n14608, QN => n8993);
   REGISTERS_reg_19_58_inst : DFF_X1 port map( D => n6659, CK => CLK, Q => 
                           n14607, QN => n8998);
   REGISTERS_reg_19_57_inst : DFF_X1 port map( D => n6658, CK => CLK, Q => 
                           n14606, QN => n9003);
   REGISTERS_reg_19_56_inst : DFF_X1 port map( D => n6657, CK => CLK, Q => 
                           n14605, QN => n9008);
   REGISTERS_reg_19_55_inst : DFF_X1 port map( D => n6656, CK => CLK, Q => 
                           n14604, QN => n9013);
   REGISTERS_reg_19_54_inst : DFF_X1 port map( D => n6655, CK => CLK, Q => 
                           n14603, QN => n9018);
   REGISTERS_reg_19_53_inst : DFF_X1 port map( D => n6654, CK => CLK, Q => 
                           n14602, QN => n9023);
   REGISTERS_reg_19_52_inst : DFF_X1 port map( D => n6653, CK => CLK, Q => 
                           n14601, QN => n9028);
   REGISTERS_reg_19_51_inst : DFF_X1 port map( D => n6652, CK => CLK, Q => 
                           n14600, QN => n9033);
   REGISTERS_reg_19_50_inst : DFF_X1 port map( D => n6651, CK => CLK, Q => 
                           n14599, QN => n9038);
   REGISTERS_reg_19_49_inst : DFF_X1 port map( D => n6650, CK => CLK, Q => 
                           n14598, QN => n9043);
   REGISTERS_reg_19_48_inst : DFF_X1 port map( D => n6649, CK => CLK, Q => 
                           n14597, QN => n9048);
   REGISTERS_reg_19_47_inst : DFF_X1 port map( D => n6648, CK => CLK, Q => 
                           n14596, QN => n9053);
   REGISTERS_reg_19_46_inst : DFF_X1 port map( D => n6647, CK => CLK, Q => 
                           n14595, QN => n9058);
   REGISTERS_reg_19_45_inst : DFF_X1 port map( D => n6646, CK => CLK, Q => 
                           n14594, QN => n9063);
   REGISTERS_reg_19_44_inst : DFF_X1 port map( D => n6645, CK => CLK, Q => 
                           n14593, QN => n9068);
   REGISTERS_reg_19_43_inst : DFF_X1 port map( D => n6644, CK => CLK, Q => 
                           n14592, QN => n9073);
   REGISTERS_reg_19_42_inst : DFF_X1 port map( D => n6643, CK => CLK, Q => 
                           n14591, QN => n9078);
   REGISTERS_reg_19_41_inst : DFF_X1 port map( D => n6642, CK => CLK, Q => 
                           n14590, QN => n9083);
   REGISTERS_reg_19_40_inst : DFF_X1 port map( D => n6641, CK => CLK, Q => 
                           n14589, QN => n9088);
   REGISTERS_reg_19_39_inst : DFF_X1 port map( D => n6640, CK => CLK, Q => 
                           n14588, QN => n9093);
   REGISTERS_reg_19_38_inst : DFF_X1 port map( D => n6639, CK => CLK, Q => 
                           n14587, QN => n9098);
   REGISTERS_reg_19_37_inst : DFF_X1 port map( D => n6638, CK => CLK, Q => 
                           n14586, QN => n9103);
   REGISTERS_reg_19_36_inst : DFF_X1 port map( D => n6637, CK => CLK, Q => 
                           n14585, QN => n9108);
   REGISTERS_reg_19_35_inst : DFF_X1 port map( D => n6636, CK => CLK, Q => 
                           n14584, QN => n9113);
   REGISTERS_reg_19_34_inst : DFF_X1 port map( D => n6635, CK => CLK, Q => 
                           n14583, QN => n9118);
   REGISTERS_reg_19_33_inst : DFF_X1 port map( D => n6634, CK => CLK, Q => 
                           n14582, QN => n9123);
   REGISTERS_reg_19_32_inst : DFF_X1 port map( D => n6633, CK => CLK, Q => 
                           n14581, QN => n9128);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n6632, CK => CLK, Q => 
                           n14580, QN => n9133);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n6631, CK => CLK, Q => 
                           n14579, QN => n9138);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n6630, CK => CLK, Q => 
                           n14578, QN => n9143);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n6629, CK => CLK, Q => 
                           n14577, QN => n9148);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n6628, CK => CLK, Q => 
                           n14576, QN => n9153);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n6627, CK => CLK, Q => 
                           n14575, QN => n9158);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n6626, CK => CLK, Q => 
                           n14574, QN => n9163);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n6625, CK => CLK, Q => 
                           n14573, QN => n9168);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n6624, CK => CLK, Q => 
                           n14572, QN => n9173);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n6623, CK => CLK, Q => 
                           n14571, QN => n9178);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n6622, CK => CLK, Q => 
                           n14570, QN => n9183);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n6621, CK => CLK, Q => 
                           n14569, QN => n9188);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n6620, CK => CLK, Q => 
                           n14568, QN => n9193);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n6619, CK => CLK, Q => 
                           n14567, QN => n9198);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n6618, CK => CLK, Q => 
                           n14566, QN => n9203);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n6617, CK => CLK, Q => 
                           n14565, QN => n9208);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n6616, CK => CLK, Q => 
                           n14564, QN => n9213);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n6615, CK => CLK, Q => 
                           n14563, QN => n9218);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n6614, CK => CLK, Q => 
                           n14562, QN => n9223);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n6613, CK => CLK, Q => 
                           n14561, QN => n9228);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n6612, CK => CLK, Q => 
                           n14560, QN => n9233);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n6611, CK => CLK, Q => 
                           n14559, QN => n9238);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n6610, CK => CLK, Q => 
                           n14558, QN => n9243);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n6609, CK => CLK, Q => 
                           n14557, QN => n9248);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n6608, CK => CLK, Q => 
                           n14556, QN => n9253);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n6607, CK => CLK, Q => 
                           n14555, QN => n9258);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n6606, CK => CLK, Q => 
                           n14554, QN => n9263);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n6605, CK => CLK, Q => 
                           n14553, QN => n9268);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n6604, CK => CLK, Q => 
                           n14552, QN => n9273);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n6603, CK => CLK, Q => 
                           n14551, QN => n9278);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n6602, CK => CLK, Q => 
                           n14550, QN => n9283);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n6601, CK => CLK, Q => 
                           n14549, QN => n9288);
   REGISTERS_reg_28_63_inst : DFF_X1 port map( D => n6088, CK => CLK, Q => 
                           n14036, QN => n9740);
   REGISTERS_reg_28_62_inst : DFF_X1 port map( D => n6087, CK => CLK, Q => 
                           n14035, QN => n9745);
   REGISTERS_reg_28_61_inst : DFF_X1 port map( D => n6086, CK => CLK, Q => 
                           n14034, QN => n9750);
   REGISTERS_reg_28_60_inst : DFF_X1 port map( D => n6085, CK => CLK, Q => 
                           n14033, QN => n9755);
   REGISTERS_reg_28_59_inst : DFF_X1 port map( D => n6084, CK => CLK, Q => 
                           n14032, QN => n9760);
   REGISTERS_reg_28_58_inst : DFF_X1 port map( D => n6083, CK => CLK, Q => 
                           n14031, QN => n9765);
   REGISTERS_reg_28_57_inst : DFF_X1 port map( D => n6082, CK => CLK, Q => 
                           n14030, QN => n9770);
   REGISTERS_reg_28_56_inst : DFF_X1 port map( D => n6081, CK => CLK, Q => 
                           n14029, QN => n9775);
   REGISTERS_reg_28_55_inst : DFF_X1 port map( D => n6080, CK => CLK, Q => 
                           n14028, QN => n9780);
   REGISTERS_reg_28_54_inst : DFF_X1 port map( D => n6079, CK => CLK, Q => 
                           n14027, QN => n9785);
   REGISTERS_reg_28_53_inst : DFF_X1 port map( D => n6078, CK => CLK, Q => 
                           n14026, QN => n9790);
   REGISTERS_reg_28_52_inst : DFF_X1 port map( D => n6077, CK => CLK, Q => 
                           n14025, QN => n9795);
   REGISTERS_reg_28_51_inst : DFF_X1 port map( D => n6076, CK => CLK, Q => 
                           n14024, QN => n9800);
   REGISTERS_reg_28_50_inst : DFF_X1 port map( D => n6075, CK => CLK, Q => 
                           n14023, QN => n9805);
   REGISTERS_reg_28_49_inst : DFF_X1 port map( D => n6074, CK => CLK, Q => 
                           n14022, QN => n9810);
   REGISTERS_reg_28_48_inst : DFF_X1 port map( D => n6073, CK => CLK, Q => 
                           n14021, QN => n9815);
   REGISTERS_reg_28_47_inst : DFF_X1 port map( D => n6072, CK => CLK, Q => 
                           n14020, QN => n9820);
   REGISTERS_reg_28_46_inst : DFF_X1 port map( D => n6071, CK => CLK, Q => 
                           n14019, QN => n9825);
   REGISTERS_reg_28_45_inst : DFF_X1 port map( D => n6070, CK => CLK, Q => 
                           n14018, QN => n9830);
   REGISTERS_reg_28_44_inst : DFF_X1 port map( D => n6069, CK => CLK, Q => 
                           n14017, QN => n9835);
   REGISTERS_reg_28_43_inst : DFF_X1 port map( D => n6068, CK => CLK, Q => 
                           n14016, QN => n9840);
   REGISTERS_reg_28_42_inst : DFF_X1 port map( D => n6067, CK => CLK, Q => 
                           n14015, QN => n9845);
   REGISTERS_reg_28_41_inst : DFF_X1 port map( D => n6066, CK => CLK, Q => 
                           n14014, QN => n9850);
   REGISTERS_reg_28_40_inst : DFF_X1 port map( D => n6065, CK => CLK, Q => 
                           n14013, QN => n9855);
   REGISTERS_reg_28_39_inst : DFF_X1 port map( D => n6064, CK => CLK, Q => 
                           n14012, QN => n9860);
   REGISTERS_reg_28_38_inst : DFF_X1 port map( D => n6063, CK => CLK, Q => 
                           n14011, QN => n9865);
   REGISTERS_reg_28_37_inst : DFF_X1 port map( D => n6062, CK => CLK, Q => 
                           n14010, QN => n9870);
   REGISTERS_reg_28_36_inst : DFF_X1 port map( D => n6061, CK => CLK, Q => 
                           n14009, QN => n9875);
   REGISTERS_reg_28_35_inst : DFF_X1 port map( D => n6060, CK => CLK, Q => 
                           n14008, QN => n9880);
   REGISTERS_reg_28_34_inst : DFF_X1 port map( D => n6059, CK => CLK, Q => 
                           n14007, QN => n9885);
   REGISTERS_reg_28_33_inst : DFF_X1 port map( D => n6058, CK => CLK, Q => 
                           n14006, QN => n9890);
   REGISTERS_reg_28_32_inst : DFF_X1 port map( D => n6057, CK => CLK, Q => 
                           n14005, QN => n9895);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n6056, CK => CLK, Q => 
                           n14004, QN => n9900);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n6055, CK => CLK, Q => 
                           n14003, QN => n9905);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n6054, CK => CLK, Q => 
                           n14002, QN => n9910);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n6053, CK => CLK, Q => 
                           n14001, QN => n9915);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n6052, CK => CLK, Q => 
                           n14000, QN => n9920);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n6051, CK => CLK, Q => 
                           n13999, QN => n9925);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n6050, CK => CLK, Q => 
                           n13998, QN => n9930);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n6049, CK => CLK, Q => 
                           n13997, QN => n9935);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n6048, CK => CLK, Q => 
                           n13996, QN => n9940);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n6047, CK => CLK, Q => 
                           n13995, QN => n9945);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n6046, CK => CLK, Q => 
                           n13994, QN => n9950);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n6045, CK => CLK, Q => 
                           n13993, QN => n9955);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n6044, CK => CLK, Q => 
                           n13992, QN => n9960);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n6043, CK => CLK, Q => 
                           n13991, QN => n9965);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n6042, CK => CLK, Q => 
                           n13990, QN => n9970);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n6041, CK => CLK, Q => 
                           n13989, QN => n9975);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n6040, CK => CLK, Q => 
                           n13988, QN => n9980);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n6039, CK => CLK, Q => 
                           n13987, QN => n9985);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n6038, CK => CLK, Q => 
                           n13986, QN => n9990);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n6037, CK => CLK, Q => 
                           n13985, QN => n9995);
   REGISTERS_reg_29_63_inst : DFF_X1 port map( D => n6024, CK => CLK, Q => 
                           n13972, QN => n8972);
   REGISTERS_reg_29_62_inst : DFF_X1 port map( D => n6023, CK => CLK, Q => 
                           n13971, QN => n8977);
   REGISTERS_reg_29_61_inst : DFF_X1 port map( D => n6022, CK => CLK, Q => 
                           n13970, QN => n8982);
   REGISTERS_reg_29_60_inst : DFF_X1 port map( D => n6021, CK => CLK, Q => 
                           n13969, QN => n8987);
   REGISTERS_reg_29_59_inst : DFF_X1 port map( D => n6020, CK => CLK, Q => 
                           n13968, QN => n8992);
   REGISTERS_reg_29_58_inst : DFF_X1 port map( D => n6019, CK => CLK, Q => 
                           n13967, QN => n8997);
   REGISTERS_reg_29_57_inst : DFF_X1 port map( D => n6018, CK => CLK, Q => 
                           n13966, QN => n9002);
   REGISTERS_reg_29_56_inst : DFF_X1 port map( D => n6017, CK => CLK, Q => 
                           n13965, QN => n9007);
   REGISTERS_reg_29_55_inst : DFF_X1 port map( D => n6016, CK => CLK, Q => 
                           n13964, QN => n9012);
   REGISTERS_reg_29_54_inst : DFF_X1 port map( D => n6015, CK => CLK, Q => 
                           n13963, QN => n9017);
   REGISTERS_reg_29_53_inst : DFF_X1 port map( D => n6014, CK => CLK, Q => 
                           n13962, QN => n9022);
   REGISTERS_reg_29_52_inst : DFF_X1 port map( D => n6013, CK => CLK, Q => 
                           n13961, QN => n9027);
   REGISTERS_reg_29_51_inst : DFF_X1 port map( D => n6012, CK => CLK, Q => 
                           n13960, QN => n9032);
   REGISTERS_reg_29_50_inst : DFF_X1 port map( D => n6011, CK => CLK, Q => 
                           n13959, QN => n9037);
   REGISTERS_reg_29_49_inst : DFF_X1 port map( D => n6010, CK => CLK, Q => 
                           n13958, QN => n9042);
   REGISTERS_reg_29_48_inst : DFF_X1 port map( D => n6009, CK => CLK, Q => 
                           n13957, QN => n9047);
   REGISTERS_reg_29_47_inst : DFF_X1 port map( D => n6008, CK => CLK, Q => 
                           n13956, QN => n9052);
   REGISTERS_reg_29_46_inst : DFF_X1 port map( D => n6007, CK => CLK, Q => 
                           n13955, QN => n9057);
   REGISTERS_reg_29_45_inst : DFF_X1 port map( D => n6006, CK => CLK, Q => 
                           n13954, QN => n9062);
   REGISTERS_reg_29_44_inst : DFF_X1 port map( D => n6005, CK => CLK, Q => 
                           n13953, QN => n9067);
   REGISTERS_reg_29_43_inst : DFF_X1 port map( D => n6004, CK => CLK, Q => 
                           n13952, QN => n9072);
   REGISTERS_reg_29_42_inst : DFF_X1 port map( D => n6003, CK => CLK, Q => 
                           n13951, QN => n9077);
   REGISTERS_reg_29_41_inst : DFF_X1 port map( D => n6002, CK => CLK, Q => 
                           n13950, QN => n9082);
   REGISTERS_reg_29_40_inst : DFF_X1 port map( D => n6001, CK => CLK, Q => 
                           n13949, QN => n9087);
   REGISTERS_reg_29_39_inst : DFF_X1 port map( D => n6000, CK => CLK, Q => 
                           n13948, QN => n9092);
   REGISTERS_reg_29_38_inst : DFF_X1 port map( D => n5999, CK => CLK, Q => 
                           n13947, QN => n9097);
   REGISTERS_reg_29_37_inst : DFF_X1 port map( D => n5998, CK => CLK, Q => 
                           n13946, QN => n9102);
   REGISTERS_reg_29_36_inst : DFF_X1 port map( D => n5997, CK => CLK, Q => 
                           n13945, QN => n9107);
   REGISTERS_reg_29_35_inst : DFF_X1 port map( D => n5996, CK => CLK, Q => 
                           n13944, QN => n9112);
   REGISTERS_reg_29_34_inst : DFF_X1 port map( D => n5995, CK => CLK, Q => 
                           n13943, QN => n9117);
   REGISTERS_reg_29_33_inst : DFF_X1 port map( D => n5994, CK => CLK, Q => 
                           n13942, QN => n9122);
   REGISTERS_reg_29_32_inst : DFF_X1 port map( D => n5993, CK => CLK, Q => 
                           n13941, QN => n9127);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n5992, CK => CLK, Q => 
                           n13940, QN => n9132);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n5991, CK => CLK, Q => 
                           n13939, QN => n9137);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n5990, CK => CLK, Q => 
                           n13938, QN => n9142);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n5989, CK => CLK, Q => 
                           n13937, QN => n9147);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n5988, CK => CLK, Q => 
                           n13936, QN => n9152);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n5987, CK => CLK, Q => 
                           n13935, QN => n9157);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n5986, CK => CLK, Q => 
                           n13934, QN => n9162);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n5985, CK => CLK, Q => 
                           n13933, QN => n9167);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n5984, CK => CLK, Q => 
                           n13932, QN => n9172);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n5983, CK => CLK, Q => 
                           n13931, QN => n9177);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n5982, CK => CLK, Q => 
                           n13930, QN => n9182);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n5981, CK => CLK, Q => 
                           n13929, QN => n9187);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n5980, CK => CLK, Q => 
                           n13928, QN => n9192);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n5979, CK => CLK, Q => 
                           n13927, QN => n9197);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n5978, CK => CLK, Q => 
                           n13926, QN => n9202);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n5977, CK => CLK, Q => 
                           n13925, QN => n9207);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n5976, CK => CLK, Q => 
                           n13924, QN => n9212);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n5975, CK => CLK, Q => 
                           n13923, QN => n9217);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n5974, CK => CLK, Q => 
                           n13922, QN => n9222);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n5973, CK => CLK, Q => 
                           n13921, QN => n9227);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n5972, CK => CLK, Q => 
                           n13920, QN => n9232);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n5971, CK => CLK, Q => 
                           n13919, QN => n9237);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n5970, CK => CLK, Q => 
                           n13918, QN => n9242);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n5969, CK => CLK, Q => 
                           n13917, QN => n9247);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n5968, CK => CLK, Q => 
                           n13916, QN => n9252);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n5967, CK => CLK, Q => 
                           n13915, QN => n9257);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n5966, CK => CLK, Q => 
                           n13914, QN => n9262);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n5965, CK => CLK, Q => 
                           n13913, QN => n9267);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n5964, CK => CLK, Q => 
                           n13912, QN => n9272);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n5963, CK => CLK, Q => 
                           n13911, QN => n9277);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n5962, CK => CLK, Q => 
                           n13910, QN => n9282);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n5961, CK => CLK, Q => 
                           n13909, QN => n9287);
   OUT2_reg_63_inst : DFF_X1 port map( D => n5895, CK => CLK, Q => n29319, QN 
                           => n10761);
   OUT2_reg_62_inst : DFF_X1 port map( D => n5893, CK => CLK, Q => n29318, QN 
                           => n10762);
   OUT2_reg_61_inst : DFF_X1 port map( D => n5891, CK => CLK, Q => n29317, QN 
                           => n10763);
   OUT2_reg_60_inst : DFF_X1 port map( D => n5889, CK => CLK, Q => n29316, QN 
                           => n10764);
   OUT2_reg_59_inst : DFF_X1 port map( D => n5887, CK => CLK, Q => n29413, QN 
                           => n10765);
   OUT2_reg_58_inst : DFF_X1 port map( D => n5885, CK => CLK, Q => n29412, QN 
                           => n10766);
   OUT2_reg_57_inst : DFF_X1 port map( D => n5883, CK => CLK, Q => n29411, QN 
                           => n10767);
   OUT2_reg_56_inst : DFF_X1 port map( D => n5881, CK => CLK, Q => n29410, QN 
                           => n10768);
   OUT2_reg_55_inst : DFF_X1 port map( D => n5879, CK => CLK, Q => n29409, QN 
                           => n10769);
   OUT2_reg_54_inst : DFF_X1 port map( D => n5877, CK => CLK, Q => n29408, QN 
                           => n10770);
   OUT2_reg_53_inst : DFF_X1 port map( D => n5875, CK => CLK, Q => n29407, QN 
                           => n10771);
   OUT2_reg_52_inst : DFF_X1 port map( D => n5873, CK => CLK, Q => n29406, QN 
                           => n10772);
   OUT2_reg_51_inst : DFF_X1 port map( D => n5871, CK => CLK, Q => n29405, QN 
                           => n10773);
   OUT2_reg_50_inst : DFF_X1 port map( D => n5869, CK => CLK, Q => n29443, QN 
                           => n10774);
   OUT2_reg_49_inst : DFF_X1 port map( D => n5867, CK => CLK, Q => n29442, QN 
                           => n10775);
   OUT2_reg_48_inst : DFF_X1 port map( D => n5865, CK => CLK, Q => n29441, QN 
                           => n10776);
   OUT2_reg_47_inst : DFF_X1 port map( D => n5863, CK => CLK, Q => n29440, QN 
                           => n10777);
   OUT2_reg_46_inst : DFF_X1 port map( D => n5861, CK => CLK, Q => n29439, QN 
                           => n10778);
   OUT2_reg_45_inst : DFF_X1 port map( D => n5859, CK => CLK, Q => n29438, QN 
                           => n10779);
   OUT2_reg_44_inst : DFF_X1 port map( D => n5857, CK => CLK, Q => n29437, QN 
                           => n10780);
   OUT2_reg_43_inst : DFF_X1 port map( D => n5855, CK => CLK, Q => n29436, QN 
                           => n10781);
   OUT2_reg_42_inst : DFF_X1 port map( D => n5853, CK => CLK, Q => n29435, QN 
                           => n10782);
   OUT2_reg_41_inst : DFF_X1 port map( D => n5851, CK => CLK, Q => n29434, QN 
                           => n10783);
   OUT2_reg_40_inst : DFF_X1 port map( D => n5849, CK => CLK, Q => n29433, QN 
                           => n10784);
   OUT2_reg_39_inst : DFF_X1 port map( D => n5847, CK => CLK, Q => n29432, QN 
                           => n10785);
   OUT2_reg_38_inst : DFF_X1 port map( D => n5845, CK => CLK, Q => n29431, QN 
                           => n10786);
   OUT2_reg_37_inst : DFF_X1 port map( D => n5843, CK => CLK, Q => n29430, QN 
                           => n10787);
   OUT2_reg_36_inst : DFF_X1 port map( D => n5841, CK => CLK, Q => n29429, QN 
                           => n10788);
   OUT2_reg_35_inst : DFF_X1 port map( D => n5839, CK => CLK, Q => n29428, QN 
                           => n10789);
   OUT2_reg_34_inst : DFF_X1 port map( D => n5837, CK => CLK, Q => n29427, QN 
                           => n10790);
   OUT2_reg_33_inst : DFF_X1 port map( D => n5835, CK => CLK, Q => n29426, QN 
                           => n10791);
   OUT2_reg_32_inst : DFF_X1 port map( D => n5833, CK => CLK, Q => n29425, QN 
                           => n10792);
   OUT2_reg_31_inst : DFF_X1 port map( D => n5831, CK => CLK, Q => n29424, QN 
                           => n10793);
   OUT2_reg_30_inst : DFF_X1 port map( D => n5829, CK => CLK, Q => n29423, QN 
                           => n10794);
   OUT2_reg_29_inst : DFF_X1 port map( D => n5827, CK => CLK, Q => n29422, QN 
                           => n10795);
   OUT2_reg_28_inst : DFF_X1 port map( D => n5825, CK => CLK, Q => n29421, QN 
                           => n10796);
   OUT2_reg_27_inst : DFF_X1 port map( D => n5823, CK => CLK, Q => n29420, QN 
                           => n10797);
   OUT2_reg_26_inst : DFF_X1 port map( D => n5821, CK => CLK, Q => n29419, QN 
                           => n10798);
   OUT2_reg_25_inst : DFF_X1 port map( D => n5819, CK => CLK, Q => n29418, QN 
                           => n10799);
   OUT2_reg_24_inst : DFF_X1 port map( D => n5817, CK => CLK, Q => n29404, QN 
                           => n10800);
   OUT2_reg_23_inst : DFF_X1 port map( D => n5815, CK => CLK, Q => n29403, QN 
                           => n10801);
   OUT2_reg_22_inst : DFF_X1 port map( D => n5813, CK => CLK, Q => n29402, QN 
                           => n10802);
   OUT2_reg_21_inst : DFF_X1 port map( D => n5811, CK => CLK, Q => n29401, QN 
                           => n10803);
   OUT2_reg_20_inst : DFF_X1 port map( D => n5809, CK => CLK, Q => n29400, QN 
                           => n10804);
   OUT2_reg_19_inst : DFF_X1 port map( D => n5807, CK => CLK, Q => n29399, QN 
                           => n10805);
   OUT2_reg_18_inst : DFF_X1 port map( D => n5805, CK => CLK, Q => n29398, QN 
                           => n10806);
   OUT2_reg_17_inst : DFF_X1 port map( D => n5803, CK => CLK, Q => n29397, QN 
                           => n10807);
   OUT2_reg_16_inst : DFF_X1 port map( D => n5801, CK => CLK, Q => n29396, QN 
                           => n10808);
   OUT2_reg_15_inst : DFF_X1 port map( D => n5799, CK => CLK, Q => n29395, QN 
                           => n10809);
   OUT2_reg_14_inst : DFF_X1 port map( D => n5797, CK => CLK, Q => n29394, QN 
                           => n10810);
   OUT2_reg_13_inst : DFF_X1 port map( D => n5795, CK => CLK, Q => n29393, QN 
                           => n10811);
   OUT2_reg_12_inst : DFF_X1 port map( D => n5793, CK => CLK, Q => n29392, QN 
                           => n10812);
   OUT2_reg_11_inst : DFF_X1 port map( D => n5791, CK => CLK, Q => n29391, QN 
                           => n10813);
   OUT2_reg_10_inst : DFF_X1 port map( D => n5789, CK => CLK, Q => n29390, QN 
                           => n10814);
   OUT2_reg_9_inst : DFF_X1 port map( D => n5787, CK => CLK, Q => n29389, QN =>
                           n10815);
   OUT2_reg_8_inst : DFF_X1 port map( D => n5785, CK => CLK, Q => n29388, QN =>
                           n10816);
   OUT2_reg_7_inst : DFF_X1 port map( D => n5783, CK => CLK, Q => n29387, QN =>
                           n10817);
   OUT2_reg_6_inst : DFF_X1 port map( D => n5781, CK => CLK, Q => n29386, QN =>
                           n10818);
   OUT2_reg_5_inst : DFF_X1 port map( D => n5779, CK => CLK, Q => n29385, QN =>
                           n10819);
   OUT2_reg_4_inst : DFF_X1 port map( D => n5777, CK => CLK, Q => n29384, QN =>
                           n10820);
   OUT2_reg_3_inst : DFF_X1 port map( D => n5775, CK => CLK, Q => n29383, QN =>
                           n10821);
   OUT2_reg_2_inst : DFF_X1 port map( D => n5773, CK => CLK, Q => n29382, QN =>
                           n10822);
   OUT2_reg_1_inst : DFF_X1 port map( D => n5771, CK => CLK, Q => n29381, QN =>
                           n10823);
   OUT2_reg_0_inst : DFF_X1 port map( D => n5769, CK => CLK, Q => n29380, QN =>
                           n10824);
   OUT1_reg_63_inst : DFF_X1 port map( D => n5768, CK => CLK, Q => n29417, QN 
                           => n10825);
   OUT1_tri_enable_reg_63_inst : DFF_X1 port map( D => n5767, CK => CLK, Q => 
                           n5258, QN => n10953);
   OUT1_reg_62_inst : DFF_X1 port map( D => n5766, CK => CLK, Q => n29416, QN 
                           => n10826);
   OUT1_tri_enable_reg_62_inst : DFF_X1 port map( D => n5765, CK => CLK, Q => 
                           n5260, QN => n10954);
   OUT1_reg_61_inst : DFF_X1 port map( D => n5764, CK => CLK, Q => n29415, QN 
                           => n10827);
   OUT1_tri_enable_reg_61_inst : DFF_X1 port map( D => n5763, CK => CLK, Q => 
                           n5262, QN => n10955);
   OUT1_reg_60_inst : DFF_X1 port map( D => n5762, CK => CLK, Q => n29414, QN 
                           => n10828);
   OUT1_tri_enable_reg_60_inst : DFF_X1 port map( D => n5761, CK => CLK, Q => 
                           n5264, QN => n10956);
   OUT1_reg_59_inst : DFF_X1 port map( D => n5760, CK => CLK, Q => n29379, QN 
                           => n10829);
   OUT1_tri_enable_reg_59_inst : DFF_X1 port map( D => n5759, CK => CLK, Q => 
                           n5266, QN => n10957);
   OUT1_reg_58_inst : DFF_X1 port map( D => n5758, CK => CLK, Q => n29378, QN 
                           => n10830);
   OUT1_tri_enable_reg_58_inst : DFF_X1 port map( D => n5757, CK => CLK, Q => 
                           n5268, QN => n10958);
   OUT1_reg_57_inst : DFF_X1 port map( D => n5756, CK => CLK, Q => n29377, QN 
                           => n10831);
   OUT1_tri_enable_reg_57_inst : DFF_X1 port map( D => n5755, CK => CLK, Q => 
                           n5270, QN => n10959);
   OUT1_reg_56_inst : DFF_X1 port map( D => n5754, CK => CLK, Q => n29376, QN 
                           => n10832);
   OUT1_tri_enable_reg_56_inst : DFF_X1 port map( D => n5753, CK => CLK, Q => 
                           n5272, QN => n10960);
   OUT1_reg_55_inst : DFF_X1 port map( D => n5752, CK => CLK, Q => n29375, QN 
                           => n10833);
   OUT1_tri_enable_reg_55_inst : DFF_X1 port map( D => n5751, CK => CLK, Q => 
                           n5274, QN => n10961);
   OUT1_reg_54_inst : DFF_X1 port map( D => n5750, CK => CLK, Q => n29374, QN 
                           => n10834);
   OUT1_tri_enable_reg_54_inst : DFF_X1 port map( D => n5749, CK => CLK, Q => 
                           n5276, QN => n10962);
   OUT1_reg_53_inst : DFF_X1 port map( D => n5748, CK => CLK, Q => n29373, QN 
                           => n10835);
   OUT1_tri_enable_reg_53_inst : DFF_X1 port map( D => n5747, CK => CLK, Q => 
                           n5278, QN => n10963);
   OUT1_reg_52_inst : DFF_X1 port map( D => n5746, CK => CLK, Q => n29372, QN 
                           => n10836);
   OUT1_tri_enable_reg_52_inst : DFF_X1 port map( D => n5745, CK => CLK, Q => 
                           n5280, QN => n10964);
   OUT1_reg_51_inst : DFF_X1 port map( D => n5744, CK => CLK, Q => n29371, QN 
                           => n10837);
   OUT1_tri_enable_reg_51_inst : DFF_X1 port map( D => n5743, CK => CLK, Q => 
                           n5282, QN => n10965);
   OUT1_reg_50_inst : DFF_X1 port map( D => n5742, CK => CLK, Q => n29370, QN 
                           => n10838);
   OUT1_tri_enable_reg_50_inst : DFF_X1 port map( D => n5741, CK => CLK, Q => 
                           n5284, QN => n10966);
   OUT1_reg_49_inst : DFF_X1 port map( D => n5740, CK => CLK, Q => n29369, QN 
                           => n10839);
   OUT1_tri_enable_reg_49_inst : DFF_X1 port map( D => n5739, CK => CLK, Q => 
                           n5286, QN => n10967);
   OUT1_reg_48_inst : DFF_X1 port map( D => n5738, CK => CLK, Q => n29368, QN 
                           => n10840);
   OUT1_tri_enable_reg_48_inst : DFF_X1 port map( D => n5737, CK => CLK, Q => 
                           n5288, QN => n10968);
   OUT1_reg_47_inst : DFF_X1 port map( D => n5736, CK => CLK, Q => n29367, QN 
                           => n10841);
   OUT1_tri_enable_reg_47_inst : DFF_X1 port map( D => n5735, CK => CLK, Q => 
                           n5290, QN => n10969);
   OUT1_reg_46_inst : DFF_X1 port map( D => n5734, CK => CLK, Q => n29366, QN 
                           => n10842);
   OUT1_tri_enable_reg_46_inst : DFF_X1 port map( D => n5733, CK => CLK, Q => 
                           n5292, QN => n10970);
   OUT1_reg_45_inst : DFF_X1 port map( D => n5732, CK => CLK, Q => n29365, QN 
                           => n10843);
   OUT1_tri_enable_reg_45_inst : DFF_X1 port map( D => n5731, CK => CLK, Q => 
                           n5294, QN => n10971);
   OUT1_reg_44_inst : DFF_X1 port map( D => n5730, CK => CLK, Q => n29364, QN 
                           => n10844);
   OUT1_tri_enable_reg_44_inst : DFF_X1 port map( D => n5729, CK => CLK, Q => 
                           n5296, QN => n10972);
   OUT1_reg_43_inst : DFF_X1 port map( D => n5728, CK => CLK, Q => n29363, QN 
                           => n10845);
   OUT1_tri_enable_reg_43_inst : DFF_X1 port map( D => n5727, CK => CLK, Q => 
                           n5298, QN => n10973);
   OUT1_reg_42_inst : DFF_X1 port map( D => n5726, CK => CLK, Q => n29362, QN 
                           => n10846);
   OUT1_tri_enable_reg_42_inst : DFF_X1 port map( D => n5725, CK => CLK, Q => 
                           n5300, QN => n10974);
   OUT1_reg_41_inst : DFF_X1 port map( D => n5724, CK => CLK, Q => n29361, QN 
                           => n10847);
   OUT1_tri_enable_reg_41_inst : DFF_X1 port map( D => n5723, CK => CLK, Q => 
                           n5302, QN => n10975);
   OUT1_reg_40_inst : DFF_X1 port map( D => n5722, CK => CLK, Q => n29360, QN 
                           => n10848);
   OUT1_tri_enable_reg_40_inst : DFF_X1 port map( D => n5721, CK => CLK, Q => 
                           n5304, QN => n10976);
   OUT1_reg_39_inst : DFF_X1 port map( D => n5720, CK => CLK, Q => n29359, QN 
                           => n10849);
   OUT1_tri_enable_reg_39_inst : DFF_X1 port map( D => n5719, CK => CLK, Q => 
                           n5306, QN => n10977);
   OUT1_reg_38_inst : DFF_X1 port map( D => n5718, CK => CLK, Q => n29358, QN 
                           => n10850);
   OUT1_tri_enable_reg_38_inst : DFF_X1 port map( D => n5717, CK => CLK, Q => 
                           n5308, QN => n10978);
   OUT1_reg_37_inst : DFF_X1 port map( D => n5716, CK => CLK, Q => n29357, QN 
                           => n10851);
   OUT1_tri_enable_reg_37_inst : DFF_X1 port map( D => n5715, CK => CLK, Q => 
                           n5310, QN => n10979);
   OUT1_reg_36_inst : DFF_X1 port map( D => n5714, CK => CLK, Q => n29356, QN 
                           => n10852);
   OUT1_tri_enable_reg_36_inst : DFF_X1 port map( D => n5713, CK => CLK, Q => 
                           n5312, QN => n10980);
   OUT1_reg_35_inst : DFF_X1 port map( D => n5712, CK => CLK, Q => n29355, QN 
                           => n10853);
   OUT1_tri_enable_reg_35_inst : DFF_X1 port map( D => n5711, CK => CLK, Q => 
                           n5314, QN => n10981);
   OUT1_reg_34_inst : DFF_X1 port map( D => n5710, CK => CLK, Q => n29354, QN 
                           => n10854);
   OUT1_tri_enable_reg_34_inst : DFF_X1 port map( D => n5709, CK => CLK, Q => 
                           n5316, QN => n10982);
   OUT1_reg_33_inst : DFF_X1 port map( D => n5708, CK => CLK, Q => n29353, QN 
                           => n10855);
   OUT1_tri_enable_reg_33_inst : DFF_X1 port map( D => n5707, CK => CLK, Q => 
                           n5318, QN => n10983);
   OUT1_reg_32_inst : DFF_X1 port map( D => n5706, CK => CLK, Q => n29352, QN 
                           => n10856);
   OUT1_tri_enable_reg_32_inst : DFF_X1 port map( D => n5705, CK => CLK, Q => 
                           n5320, QN => n10984);
   OUT1_reg_31_inst : DFF_X1 port map( D => n5704, CK => CLK, Q => n29351, QN 
                           => n10857);
   OUT1_tri_enable_reg_31_inst : DFF_X1 port map( D => n5703, CK => CLK, Q => 
                           n5322, QN => n10985);
   OUT1_reg_30_inst : DFF_X1 port map( D => n5702, CK => CLK, Q => n29350, QN 
                           => n10858);
   OUT1_tri_enable_reg_30_inst : DFF_X1 port map( D => n5701, CK => CLK, Q => 
                           n5324, QN => n10986);
   OUT1_reg_29_inst : DFF_X1 port map( D => n5700, CK => CLK, Q => n29349, QN 
                           => n10859);
   OUT1_tri_enable_reg_29_inst : DFF_X1 port map( D => n5699, CK => CLK, Q => 
                           n5326, QN => n10987);
   OUT1_reg_28_inst : DFF_X1 port map( D => n5698, CK => CLK, Q => n29348, QN 
                           => n10860);
   OUT1_tri_enable_reg_28_inst : DFF_X1 port map( D => n5697, CK => CLK, Q => 
                           n5328, QN => n10988);
   OUT1_reg_27_inst : DFF_X1 port map( D => n5696, CK => CLK, Q => n29347, QN 
                           => n10861);
   OUT1_tri_enable_reg_27_inst : DFF_X1 port map( D => n5695, CK => CLK, Q => 
                           n5330, QN => n10989);
   OUT1_reg_26_inst : DFF_X1 port map( D => n5694, CK => CLK, Q => n29346, QN 
                           => n10862);
   OUT1_tri_enable_reg_26_inst : DFF_X1 port map( D => n5693, CK => CLK, Q => 
                           n5332, QN => n10990);
   OUT1_reg_25_inst : DFF_X1 port map( D => n5692, CK => CLK, Q => n29345, QN 
                           => n10863);
   OUT1_tri_enable_reg_25_inst : DFF_X1 port map( D => n5691, CK => CLK, Q => 
                           n5334, QN => n10991);
   OUT1_reg_24_inst : DFF_X1 port map( D => n5690, CK => CLK, Q => n29344, QN 
                           => n10864);
   OUT1_tri_enable_reg_24_inst : DFF_X1 port map( D => n5689, CK => CLK, Q => 
                           n5336, QN => n10992);
   OUT1_reg_23_inst : DFF_X1 port map( D => n5688, CK => CLK, Q => n29343, QN 
                           => n10865);
   OUT1_tri_enable_reg_23_inst : DFF_X1 port map( D => n5687, CK => CLK, Q => 
                           n5338, QN => n10993);
   OUT1_reg_22_inst : DFF_X1 port map( D => n5686, CK => CLK, Q => n29342, QN 
                           => n10866);
   OUT1_tri_enable_reg_22_inst : DFF_X1 port map( D => n5685, CK => CLK, Q => 
                           n5340, QN => n10994);
   OUT1_reg_21_inst : DFF_X1 port map( D => n5684, CK => CLK, Q => n29341, QN 
                           => n10867);
   OUT1_tri_enable_reg_21_inst : DFF_X1 port map( D => n5683, CK => CLK, Q => 
                           n5342, QN => n10995);
   OUT1_reg_20_inst : DFF_X1 port map( D => n5682, CK => CLK, Q => n29340, QN 
                           => n10868);
   OUT1_tri_enable_reg_20_inst : DFF_X1 port map( D => n5681, CK => CLK, Q => 
                           n5344, QN => n10996);
   OUT1_reg_19_inst : DFF_X1 port map( D => n5680, CK => CLK, Q => n29339, QN 
                           => n10869);
   OUT1_tri_enable_reg_19_inst : DFF_X1 port map( D => n5679, CK => CLK, Q => 
                           n5346, QN => n10997);
   OUT1_reg_18_inst : DFF_X1 port map( D => n5678, CK => CLK, Q => n29338, QN 
                           => n10870);
   OUT1_tri_enable_reg_18_inst : DFF_X1 port map( D => n5677, CK => CLK, Q => 
                           n5348, QN => n10998);
   OUT1_reg_17_inst : DFF_X1 port map( D => n5676, CK => CLK, Q => n29337, QN 
                           => n10871);
   OUT1_tri_enable_reg_17_inst : DFF_X1 port map( D => n5675, CK => CLK, Q => 
                           n5350, QN => n10999);
   OUT1_reg_16_inst : DFF_X1 port map( D => n5674, CK => CLK, Q => n29336, QN 
                           => n10872);
   OUT1_tri_enable_reg_16_inst : DFF_X1 port map( D => n5673, CK => CLK, Q => 
                           n5352, QN => n11000);
   OUT1_reg_15_inst : DFF_X1 port map( D => n5672, CK => CLK, Q => n29335, QN 
                           => n10873);
   OUT1_tri_enable_reg_15_inst : DFF_X1 port map( D => n5671, CK => CLK, Q => 
                           n5354, QN => n11001);
   OUT1_reg_14_inst : DFF_X1 port map( D => n5670, CK => CLK, Q => n29334, QN 
                           => n10874);
   OUT1_tri_enable_reg_14_inst : DFF_X1 port map( D => n5669, CK => CLK, Q => 
                           n5356, QN => n11002);
   OUT1_reg_13_inst : DFF_X1 port map( D => n5668, CK => CLK, Q => n29333, QN 
                           => n10875);
   OUT1_tri_enable_reg_13_inst : DFF_X1 port map( D => n5667, CK => CLK, Q => 
                           n5358, QN => n11003);
   OUT1_reg_12_inst : DFF_X1 port map( D => n5666, CK => CLK, Q => n29332, QN 
                           => n10876);
   OUT1_tri_enable_reg_12_inst : DFF_X1 port map( D => n5665, CK => CLK, Q => 
                           n5360, QN => n11004);
   OUT1_reg_11_inst : DFF_X1 port map( D => n5664, CK => CLK, Q => n29331, QN 
                           => n10877);
   OUT1_tri_enable_reg_11_inst : DFF_X1 port map( D => n5663, CK => CLK, Q => 
                           n5362, QN => n11005);
   OUT1_reg_10_inst : DFF_X1 port map( D => n5662, CK => CLK, Q => n29330, QN 
                           => n10878);
   OUT1_tri_enable_reg_10_inst : DFF_X1 port map( D => n5661, CK => CLK, Q => 
                           n5364, QN => n11006);
   OUT1_reg_9_inst : DFF_X1 port map( D => n5660, CK => CLK, Q => n29329, QN =>
                           n10879);
   OUT1_tri_enable_reg_9_inst : DFF_X1 port map( D => n5659, CK => CLK, Q => 
                           n5366, QN => n11007);
   OUT1_reg_8_inst : DFF_X1 port map( D => n5658, CK => CLK, Q => n29328, QN =>
                           n10880);
   OUT1_tri_enable_reg_8_inst : DFF_X1 port map( D => n5657, CK => CLK, Q => 
                           n5368, QN => n11008);
   OUT1_reg_7_inst : DFF_X1 port map( D => n5656, CK => CLK, Q => n29327, QN =>
                           n10881);
   OUT1_tri_enable_reg_7_inst : DFF_X1 port map( D => n5655, CK => CLK, Q => 
                           n5370, QN => n11009);
   OUT1_reg_6_inst : DFF_X1 port map( D => n5654, CK => CLK, Q => n29326, QN =>
                           n10882);
   OUT1_tri_enable_reg_6_inst : DFF_X1 port map( D => n5653, CK => CLK, Q => 
                           n5372, QN => n11010);
   OUT1_reg_5_inst : DFF_X1 port map( D => n5652, CK => CLK, Q => n29325, QN =>
                           n10883);
   OUT1_tri_enable_reg_5_inst : DFF_X1 port map( D => n5651, CK => CLK, Q => 
                           n5374, QN => n11011);
   OUT1_reg_4_inst : DFF_X1 port map( D => n5650, CK => CLK, Q => n29324, QN =>
                           n10884);
   OUT1_tri_enable_reg_4_inst : DFF_X1 port map( D => n5649, CK => CLK, Q => 
                           n5376, QN => n11012);
   OUT1_reg_3_inst : DFF_X1 port map( D => n5648, CK => CLK, Q => n29323, QN =>
                           n10885);
   OUT1_tri_enable_reg_3_inst : DFF_X1 port map( D => n5647, CK => CLK, Q => 
                           n5378, QN => n11013);
   OUT1_reg_2_inst : DFF_X1 port map( D => n5646, CK => CLK, Q => n29322, QN =>
                           n10886);
   OUT1_tri_enable_reg_2_inst : DFF_X1 port map( D => n5645, CK => CLK, Q => 
                           n5380, QN => n11014);
   OUT1_reg_1_inst : DFF_X1 port map( D => n5644, CK => CLK, Q => n29321, QN =>
                           n10887);
   OUT1_tri_enable_reg_1_inst : DFF_X1 port map( D => n5643, CK => CLK, Q => 
                           n5382, QN => n11015);
   OUT1_reg_0_inst : DFF_X1 port map( D => n5642, CK => CLK, Q => n29320, QN =>
                           n10888);
   OUT1_tri_enable_reg_0_inst : DFF_X1 port map( D => n5641, CK => CLK, Q => 
                           n5384, QN => n11016);
   REGISTERS_reg_24_63_inst : DFF_X1 port map( D => n6344, CK => CLK, Q => 
                           n29507, QN => n18192);
   REGISTERS_reg_24_62_inst : DFF_X1 port map( D => n6343, CK => CLK, Q => 
                           n29506, QN => n18194);
   REGISTERS_reg_24_61_inst : DFF_X1 port map( D => n6342, CK => CLK, Q => 
                           n29505, QN => n18195);
   REGISTERS_reg_24_60_inst : DFF_X1 port map( D => n6341, CK => CLK, Q => 
                           n29504, QN => n18196);
   REGISTERS_reg_23_63_inst : DFF_X1 port map( D => n6408, CK => CLK, Q => 
                           n29763, QN => n18126);
   REGISTERS_reg_23_62_inst : DFF_X1 port map( D => n6407, CK => CLK, Q => 
                           n29762, QN => n18128);
   REGISTERS_reg_23_61_inst : DFF_X1 port map( D => n6406, CK => CLK, Q => 
                           n29761, QN => n18129);
   REGISTERS_reg_23_60_inst : DFF_X1 port map( D => n6405, CK => CLK, Q => 
                           n29760, QN => n18130);
   REGISTERS_reg_25_63_inst : DFF_X1 port map( D => n6280, CK => CLK, Q => 
                           n29699, QN => n18259);
   REGISTERS_reg_25_62_inst : DFF_X1 port map( D => n6279, CK => CLK, Q => 
                           n29698, QN => n18261);
   REGISTERS_reg_25_61_inst : DFF_X1 port map( D => n6278, CK => CLK, Q => 
                           n29697, QN => n18262);
   REGISTERS_reg_25_60_inst : DFF_X1 port map( D => n6277, CK => CLK, Q => 
                           n29696, QN => n18263);
   REGISTERS_reg_22_63_inst : DFF_X1 port map( D => n6472, CK => CLK, Q => 
                           n29571, QN => n18059);
   REGISTERS_reg_22_62_inst : DFF_X1 port map( D => n6471, CK => CLK, Q => 
                           n29570, QN => n18061);
   REGISTERS_reg_22_61_inst : DFF_X1 port map( D => n6470, CK => CLK, Q => 
                           n29569, QN => n18062);
   REGISTERS_reg_22_60_inst : DFF_X1 port map( D => n6469, CK => CLK, Q => 
                           n29568, QN => n18063);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n6356, CK => CLK, Q => 
                           n29711, QN => n18179);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n6355, CK => CLK, Q => 
                           n29710, QN => n18180);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n6354, CK => CLK, Q => 
                           n29709, QN => n18181);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n6353, CK => CLK, Q => 
                           n29708, QN => n18182);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n6352, CK => CLK, Q => 
                           n29707, QN => n18183);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n6351, CK => CLK, Q => 
                           n29706, QN => n18184);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n6350, CK => CLK, Q => 
                           n29705, QN => n18185);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n6349, CK => CLK, Q => 
                           n29704, QN => n18186);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n6348, CK => CLK, Q => 
                           n29703, QN => n18187);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n6347, CK => CLK, Q => 
                           n29702, QN => n18188);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n6346, CK => CLK, Q => 
                           n29701, QN => n18189);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n6345, CK => CLK, Q => 
                           n29700, QN => n18190);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n6420, CK => CLK, Q => 
                           n29519, QN => n18112);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n6419, CK => CLK, Q => 
                           n29518, QN => n18113);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n6418, CK => CLK, Q => 
                           n29517, QN => n18114);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n6417, CK => CLK, Q => 
                           n29516, QN => n18115);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n6416, CK => CLK, Q => 
                           n29515, QN => n18116);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n6415, CK => CLK, Q => 
                           n29514, QN => n18117);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n6414, CK => CLK, Q => 
                           n29513, QN => n18118);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n6413, CK => CLK, Q => 
                           n29512, QN => n18119);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n6412, CK => CLK, Q => 
                           n29511, QN => n18120);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n6411, CK => CLK, Q => 
                           n29510, QN => n18121);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n6410, CK => CLK, Q => 
                           n29509, QN => n18122);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n6409, CK => CLK, Q => 
                           n29508, QN => n18123);
   REGISTERS_reg_23_59_inst : DFF_X1 port map( D => n6404, CK => CLK, Q => 
                           n29759, QN => n18131);
   REGISTERS_reg_23_58_inst : DFF_X1 port map( D => n6403, CK => CLK, Q => 
                           n29758, QN => n18132);
   REGISTERS_reg_23_57_inst : DFF_X1 port map( D => n6402, CK => CLK, Q => 
                           n29757, QN => n18133);
   REGISTERS_reg_23_56_inst : DFF_X1 port map( D => n6401, CK => CLK, Q => 
                           n29756, QN => n18134);
   REGISTERS_reg_23_55_inst : DFF_X1 port map( D => n6400, CK => CLK, Q => 
                           n29755, QN => n18135);
   REGISTERS_reg_23_54_inst : DFF_X1 port map( D => n6399, CK => CLK, Q => 
                           n29754, QN => n18136);
   REGISTERS_reg_23_53_inst : DFF_X1 port map( D => n6398, CK => CLK, Q => 
                           n29753, QN => n18137);
   REGISTERS_reg_23_52_inst : DFF_X1 port map( D => n6397, CK => CLK, Q => 
                           n29752, QN => n18138);
   REGISTERS_reg_23_51_inst : DFF_X1 port map( D => n6396, CK => CLK, Q => 
                           n29751, QN => n18139);
   REGISTERS_reg_23_50_inst : DFF_X1 port map( D => n6395, CK => CLK, Q => 
                           n29750, QN => n18140);
   REGISTERS_reg_23_49_inst : DFF_X1 port map( D => n6394, CK => CLK, Q => 
                           n29749, QN => n18141);
   REGISTERS_reg_23_48_inst : DFF_X1 port map( D => n6393, CK => CLK, Q => 
                           n29748, QN => n18142);
   REGISTERS_reg_23_47_inst : DFF_X1 port map( D => n6392, CK => CLK, Q => 
                           n29747, QN => n18143);
   REGISTERS_reg_23_46_inst : DFF_X1 port map( D => n6391, CK => CLK, Q => 
                           n29746, QN => n18144);
   REGISTERS_reg_23_45_inst : DFF_X1 port map( D => n6390, CK => CLK, Q => 
                           n29745, QN => n18145);
   REGISTERS_reg_23_44_inst : DFF_X1 port map( D => n6389, CK => CLK, Q => 
                           n29744, QN => n18146);
   REGISTERS_reg_23_43_inst : DFF_X1 port map( D => n6388, CK => CLK, Q => 
                           n29743, QN => n18147);
   REGISTERS_reg_23_42_inst : DFF_X1 port map( D => n6387, CK => CLK, Q => 
                           n29742, QN => n18148);
   REGISTERS_reg_23_41_inst : DFF_X1 port map( D => n6386, CK => CLK, Q => 
                           n29741, QN => n18149);
   REGISTERS_reg_23_40_inst : DFF_X1 port map( D => n6385, CK => CLK, Q => 
                           n29740, QN => n18150);
   REGISTERS_reg_23_39_inst : DFF_X1 port map( D => n6384, CK => CLK, Q => 
                           n29739, QN => n18151);
   REGISTERS_reg_23_38_inst : DFF_X1 port map( D => n6383, CK => CLK, Q => 
                           n29738, QN => n18152);
   REGISTERS_reg_23_37_inst : DFF_X1 port map( D => n6382, CK => CLK, Q => 
                           n29737, QN => n18153);
   REGISTERS_reg_23_36_inst : DFF_X1 port map( D => n6381, CK => CLK, Q => 
                           n29736, QN => n18154);
   REGISTERS_reg_23_35_inst : DFF_X1 port map( D => n6380, CK => CLK, Q => 
                           n29735, QN => n18155);
   REGISTERS_reg_23_34_inst : DFF_X1 port map( D => n6379, CK => CLK, Q => 
                           n29734, QN => n18156);
   REGISTERS_reg_23_33_inst : DFF_X1 port map( D => n6378, CK => CLK, Q => 
                           n29733, QN => n18157);
   REGISTERS_reg_23_32_inst : DFF_X1 port map( D => n6377, CK => CLK, Q => 
                           n29732, QN => n18158);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n6376, CK => CLK, Q => 
                           n29731, QN => n18159);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n6375, CK => CLK, Q => 
                           n29730, QN => n18160);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n6374, CK => CLK, Q => 
                           n29729, QN => n18161);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n6373, CK => CLK, Q => 
                           n29728, QN => n18162);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n6372, CK => CLK, Q => 
                           n29727, QN => n18163);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n6371, CK => CLK, Q => 
                           n29726, QN => n18164);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n6370, CK => CLK, Q => 
                           n29725, QN => n18165);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n6369, CK => CLK, Q => 
                           n29724, QN => n18166);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n6368, CK => CLK, Q => 
                           n29723, QN => n18167);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n6367, CK => CLK, Q => 
                           n29722, QN => n18168);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n6366, CK => CLK, Q => 
                           n29721, QN => n18169);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n6365, CK => CLK, Q => 
                           n29720, QN => n18170);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n6364, CK => CLK, Q => 
                           n29719, QN => n18171);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n6363, CK => CLK, Q => 
                           n29718, QN => n18172);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n6362, CK => CLK, Q => 
                           n29717, QN => n18173);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n6361, CK => CLK, Q => 
                           n29716, QN => n18174);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n6360, CK => CLK, Q => 
                           n29715, QN => n18175);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n6359, CK => CLK, Q => 
                           n29714, QN => n18176);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n6358, CK => CLK, Q => 
                           n29713, QN => n18177);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n6357, CK => CLK, Q => 
                           n29712, QN => n18178);
   REGISTERS_reg_22_59_inst : DFF_X1 port map( D => n6468, CK => CLK, Q => 
                           n29567, QN => n18064);
   REGISTERS_reg_22_58_inst : DFF_X1 port map( D => n6467, CK => CLK, Q => 
                           n29566, QN => n18065);
   REGISTERS_reg_22_57_inst : DFF_X1 port map( D => n6466, CK => CLK, Q => 
                           n29565, QN => n18066);
   REGISTERS_reg_22_56_inst : DFF_X1 port map( D => n6465, CK => CLK, Q => 
                           n29564, QN => n18067);
   REGISTERS_reg_22_55_inst : DFF_X1 port map( D => n6464, CK => CLK, Q => 
                           n29563, QN => n18068);
   REGISTERS_reg_22_54_inst : DFF_X1 port map( D => n6463, CK => CLK, Q => 
                           n29562, QN => n18069);
   REGISTERS_reg_22_53_inst : DFF_X1 port map( D => n6462, CK => CLK, Q => 
                           n29561, QN => n18070);
   REGISTERS_reg_22_52_inst : DFF_X1 port map( D => n6461, CK => CLK, Q => 
                           n29560, QN => n18071);
   REGISTERS_reg_22_51_inst : DFF_X1 port map( D => n6460, CK => CLK, Q => 
                           n29559, QN => n18072);
   REGISTERS_reg_22_50_inst : DFF_X1 port map( D => n6459, CK => CLK, Q => 
                           n29558, QN => n18073);
   REGISTERS_reg_22_49_inst : DFF_X1 port map( D => n6458, CK => CLK, Q => 
                           n29557, QN => n18074);
   REGISTERS_reg_22_48_inst : DFF_X1 port map( D => n6457, CK => CLK, Q => 
                           n29556, QN => n18075);
   REGISTERS_reg_22_47_inst : DFF_X1 port map( D => n6456, CK => CLK, Q => 
                           n29555, QN => n18076);
   REGISTERS_reg_22_46_inst : DFF_X1 port map( D => n6455, CK => CLK, Q => 
                           n29554, QN => n18077);
   REGISTERS_reg_22_45_inst : DFF_X1 port map( D => n6454, CK => CLK, Q => 
                           n29553, QN => n18078);
   REGISTERS_reg_22_44_inst : DFF_X1 port map( D => n6453, CK => CLK, Q => 
                           n29552, QN => n18079);
   REGISTERS_reg_22_43_inst : DFF_X1 port map( D => n6452, CK => CLK, Q => 
                           n29551, QN => n18080);
   REGISTERS_reg_22_42_inst : DFF_X1 port map( D => n6451, CK => CLK, Q => 
                           n29550, QN => n18081);
   REGISTERS_reg_22_41_inst : DFF_X1 port map( D => n6450, CK => CLK, Q => 
                           n29549, QN => n18082);
   REGISTERS_reg_22_40_inst : DFF_X1 port map( D => n6449, CK => CLK, Q => 
                           n29548, QN => n18083);
   REGISTERS_reg_22_39_inst : DFF_X1 port map( D => n6448, CK => CLK, Q => 
                           n29547, QN => n18084);
   REGISTERS_reg_22_38_inst : DFF_X1 port map( D => n6447, CK => CLK, Q => 
                           n29546, QN => n18085);
   REGISTERS_reg_22_37_inst : DFF_X1 port map( D => n6446, CK => CLK, Q => 
                           n29545, QN => n18086);
   REGISTERS_reg_22_36_inst : DFF_X1 port map( D => n6445, CK => CLK, Q => 
                           n29544, QN => n18087);
   REGISTERS_reg_22_35_inst : DFF_X1 port map( D => n6444, CK => CLK, Q => 
                           n29543, QN => n18088);
   REGISTERS_reg_22_34_inst : DFF_X1 port map( D => n6443, CK => CLK, Q => 
                           n29542, QN => n18089);
   REGISTERS_reg_22_33_inst : DFF_X1 port map( D => n6442, CK => CLK, Q => 
                           n29541, QN => n18090);
   REGISTERS_reg_22_32_inst : DFF_X1 port map( D => n6441, CK => CLK, Q => 
                           n29540, QN => n18091);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n6440, CK => CLK, Q => 
                           n29539, QN => n18092);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n6439, CK => CLK, Q => 
                           n29538, QN => n18093);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n6438, CK => CLK, Q => 
                           n29537, QN => n18094);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n6437, CK => CLK, Q => 
                           n29536, QN => n18095);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n6436, CK => CLK, Q => 
                           n29535, QN => n18096);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n6435, CK => CLK, Q => 
                           n29534, QN => n18097);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n6434, CK => CLK, Q => 
                           n29533, QN => n18098);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n6433, CK => CLK, Q => 
                           n29532, QN => n18099);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n6432, CK => CLK, Q => 
                           n29531, QN => n18100);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n6431, CK => CLK, Q => 
                           n29530, QN => n18101);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n6430, CK => CLK, Q => 
                           n29529, QN => n18102);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n6429, CK => CLK, Q => 
                           n29528, QN => n18103);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n6428, CK => CLK, Q => 
                           n29527, QN => n18104);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n6427, CK => CLK, Q => 
                           n29526, QN => n18105);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n6426, CK => CLK, Q => 
                           n29525, QN => n18106);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n6425, CK => CLK, Q => 
                           n29524, QN => n18107);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n6424, CK => CLK, Q => 
                           n29523, QN => n18108);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n6423, CK => CLK, Q => 
                           n29522, QN => n18109);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n6422, CK => CLK, Q => 
                           n29521, QN => n18110);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n6421, CK => CLK, Q => 
                           n29520, QN => n18111);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n6228, CK => CLK, Q => 
                           n29647, QN => n18312);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n6227, CK => CLK, Q => 
                           n29646, QN => n18313);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n6226, CK => CLK, Q => 
                           n29645, QN => n18314);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n6225, CK => CLK, Q => 
                           n29644, QN => n18315);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n6224, CK => CLK, Q => 
                           n29643, QN => n18316);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n6223, CK => CLK, Q => 
                           n29642, QN => n18317);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n6222, CK => CLK, Q => 
                           n29641, QN => n18318);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n6221, CK => CLK, Q => 
                           n29640, QN => n18319);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n6220, CK => CLK, Q => 
                           n29639, QN => n18320);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n6219, CK => CLK, Q => 
                           n29638, QN => n18321);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n6218, CK => CLK, Q => 
                           n29637, QN => n18322);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n6217, CK => CLK, Q => 
                           n29636, QN => n18323);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n6292, CK => CLK, Q => 
                           n29455, QN => n18245);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n6291, CK => CLK, Q => 
                           n29454, QN => n18246);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n6290, CK => CLK, Q => 
                           n29453, QN => n18247);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n6289, CK => CLK, Q => 
                           n29452, QN => n18248);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n6288, CK => CLK, Q => 
                           n29451, QN => n18249);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n6287, CK => CLK, Q => 
                           n29450, QN => n18250);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n6286, CK => CLK, Q => 
                           n29449, QN => n18251);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n6285, CK => CLK, Q => 
                           n29448, QN => n18252);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n6284, CK => CLK, Q => 
                           n29447, QN => n18253);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n6283, CK => CLK, Q => 
                           n29446, QN => n18254);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n6282, CK => CLK, Q => 
                           n29445, QN => n18255);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n6281, CK => CLK, Q => 
                           n29444, QN => n18256);
   REGISTERS_reg_25_59_inst : DFF_X1 port map( D => n6276, CK => CLK, Q => 
                           n29695, QN => n18264);
   REGISTERS_reg_25_58_inst : DFF_X1 port map( D => n6275, CK => CLK, Q => 
                           n29694, QN => n18265);
   REGISTERS_reg_25_57_inst : DFF_X1 port map( D => n6274, CK => CLK, Q => 
                           n29693, QN => n18266);
   REGISTERS_reg_25_56_inst : DFF_X1 port map( D => n6273, CK => CLK, Q => 
                           n29692, QN => n18267);
   REGISTERS_reg_25_55_inst : DFF_X1 port map( D => n6272, CK => CLK, Q => 
                           n29691, QN => n18268);
   REGISTERS_reg_25_54_inst : DFF_X1 port map( D => n6271, CK => CLK, Q => 
                           n29690, QN => n18269);
   REGISTERS_reg_25_53_inst : DFF_X1 port map( D => n6270, CK => CLK, Q => 
                           n29689, QN => n18270);
   REGISTERS_reg_25_52_inst : DFF_X1 port map( D => n6269, CK => CLK, Q => 
                           n29688, QN => n18271);
   REGISTERS_reg_25_51_inst : DFF_X1 port map( D => n6268, CK => CLK, Q => 
                           n29687, QN => n18272);
   REGISTERS_reg_25_50_inst : DFF_X1 port map( D => n6267, CK => CLK, Q => 
                           n29686, QN => n18273);
   REGISTERS_reg_25_49_inst : DFF_X1 port map( D => n6266, CK => CLK, Q => 
                           n29685, QN => n18274);
   REGISTERS_reg_25_48_inst : DFF_X1 port map( D => n6265, CK => CLK, Q => 
                           n29684, QN => n18275);
   REGISTERS_reg_25_47_inst : DFF_X1 port map( D => n6264, CK => CLK, Q => 
                           n29683, QN => n18276);
   REGISTERS_reg_25_46_inst : DFF_X1 port map( D => n6263, CK => CLK, Q => 
                           n29682, QN => n18277);
   REGISTERS_reg_25_45_inst : DFF_X1 port map( D => n6262, CK => CLK, Q => 
                           n29681, QN => n18278);
   REGISTERS_reg_25_44_inst : DFF_X1 port map( D => n6261, CK => CLK, Q => 
                           n29680, QN => n18279);
   REGISTERS_reg_25_43_inst : DFF_X1 port map( D => n6260, CK => CLK, Q => 
                           n29679, QN => n18280);
   REGISTERS_reg_25_42_inst : DFF_X1 port map( D => n6259, CK => CLK, Q => 
                           n29678, QN => n18281);
   REGISTERS_reg_25_41_inst : DFF_X1 port map( D => n6258, CK => CLK, Q => 
                           n29677, QN => n18282);
   REGISTERS_reg_25_40_inst : DFF_X1 port map( D => n6257, CK => CLK, Q => 
                           n29676, QN => n18283);
   REGISTERS_reg_25_39_inst : DFF_X1 port map( D => n6256, CK => CLK, Q => 
                           n29675, QN => n18284);
   REGISTERS_reg_25_38_inst : DFF_X1 port map( D => n6255, CK => CLK, Q => 
                           n29674, QN => n18285);
   REGISTERS_reg_24_59_inst : DFF_X1 port map( D => n6340, CK => CLK, Q => 
                           n29503, QN => n18197);
   REGISTERS_reg_24_58_inst : DFF_X1 port map( D => n6339, CK => CLK, Q => 
                           n29502, QN => n18198);
   REGISTERS_reg_24_57_inst : DFF_X1 port map( D => n6338, CK => CLK, Q => 
                           n29501, QN => n18199);
   REGISTERS_reg_24_56_inst : DFF_X1 port map( D => n6337, CK => CLK, Q => 
                           n29500, QN => n18200);
   REGISTERS_reg_24_55_inst : DFF_X1 port map( D => n6336, CK => CLK, Q => 
                           n29499, QN => n18201);
   REGISTERS_reg_24_54_inst : DFF_X1 port map( D => n6335, CK => CLK, Q => 
                           n29498, QN => n18202);
   REGISTERS_reg_24_53_inst : DFF_X1 port map( D => n6334, CK => CLK, Q => 
                           n29497, QN => n18203);
   REGISTERS_reg_24_52_inst : DFF_X1 port map( D => n6333, CK => CLK, Q => 
                           n29496, QN => n18204);
   REGISTERS_reg_24_51_inst : DFF_X1 port map( D => n6332, CK => CLK, Q => 
                           n29495, QN => n18205);
   REGISTERS_reg_24_50_inst : DFF_X1 port map( D => n6331, CK => CLK, Q => 
                           n29494, QN => n18206);
   REGISTERS_reg_24_49_inst : DFF_X1 port map( D => n6330, CK => CLK, Q => 
                           n29493, QN => n18207);
   REGISTERS_reg_24_48_inst : DFF_X1 port map( D => n6329, CK => CLK, Q => 
                           n29492, QN => n18208);
   REGISTERS_reg_24_47_inst : DFF_X1 port map( D => n6328, CK => CLK, Q => 
                           n29491, QN => n18209);
   REGISTERS_reg_24_46_inst : DFF_X1 port map( D => n6327, CK => CLK, Q => 
                           n29490, QN => n18210);
   REGISTERS_reg_24_45_inst : DFF_X1 port map( D => n6326, CK => CLK, Q => 
                           n29489, QN => n18211);
   REGISTERS_reg_24_44_inst : DFF_X1 port map( D => n6325, CK => CLK, Q => 
                           n29488, QN => n18212);
   REGISTERS_reg_24_43_inst : DFF_X1 port map( D => n6324, CK => CLK, Q => 
                           n29487, QN => n18213);
   REGISTERS_reg_24_42_inst : DFF_X1 port map( D => n6323, CK => CLK, Q => 
                           n29486, QN => n18214);
   REGISTERS_reg_24_41_inst : DFF_X1 port map( D => n6322, CK => CLK, Q => 
                           n29485, QN => n18215);
   REGISTERS_reg_24_40_inst : DFF_X1 port map( D => n6321, CK => CLK, Q => 
                           n29484, QN => n18216);
   REGISTERS_reg_24_39_inst : DFF_X1 port map( D => n6320, CK => CLK, Q => 
                           n29483, QN => n18217);
   REGISTERS_reg_24_38_inst : DFF_X1 port map( D => n6319, CK => CLK, Q => 
                           n29482, QN => n18218);
   REGISTERS_reg_25_37_inst : DFF_X1 port map( D => n6254, CK => CLK, Q => 
                           n29673, QN => n18286);
   REGISTERS_reg_25_36_inst : DFF_X1 port map( D => n6253, CK => CLK, Q => 
                           n29672, QN => n18287);
   REGISTERS_reg_25_35_inst : DFF_X1 port map( D => n6252, CK => CLK, Q => 
                           n29671, QN => n18288);
   REGISTERS_reg_25_34_inst : DFF_X1 port map( D => n6251, CK => CLK, Q => 
                           n29670, QN => n18289);
   REGISTERS_reg_25_33_inst : DFF_X1 port map( D => n6250, CK => CLK, Q => 
                           n29669, QN => n18290);
   REGISTERS_reg_25_32_inst : DFF_X1 port map( D => n6249, CK => CLK, Q => 
                           n29668, QN => n18291);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n6248, CK => CLK, Q => 
                           n29667, QN => n18292);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n6247, CK => CLK, Q => 
                           n29666, QN => n18293);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n6246, CK => CLK, Q => 
                           n29665, QN => n18294);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n6245, CK => CLK, Q => 
                           n29664, QN => n18295);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n6244, CK => CLK, Q => 
                           n29663, QN => n18296);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n6243, CK => CLK, Q => 
                           n29662, QN => n18297);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n6242, CK => CLK, Q => 
                           n29661, QN => n18298);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n6241, CK => CLK, Q => 
                           n29660, QN => n18299);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n6240, CK => CLK, Q => 
                           n29659, QN => n18300);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n6239, CK => CLK, Q => 
                           n29658, QN => n18301);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n6238, CK => CLK, Q => 
                           n29657, QN => n18302);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n6237, CK => CLK, Q => 
                           n29656, QN => n18303);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n6236, CK => CLK, Q => 
                           n29655, QN => n18304);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n6235, CK => CLK, Q => 
                           n29654, QN => n18305);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n6234, CK => CLK, Q => 
                           n29653, QN => n18306);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n6233, CK => CLK, Q => 
                           n29652, QN => n18307);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n6232, CK => CLK, Q => 
                           n29651, QN => n18308);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n6231, CK => CLK, Q => 
                           n29650, QN => n18309);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n6230, CK => CLK, Q => 
                           n29649, QN => n18310);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n6229, CK => CLK, Q => 
                           n29648, QN => n18311);
   REGISTERS_reg_24_37_inst : DFF_X1 port map( D => n6318, CK => CLK, Q => 
                           n29481, QN => n18219);
   REGISTERS_reg_24_36_inst : DFF_X1 port map( D => n6317, CK => CLK, Q => 
                           n29480, QN => n18220);
   REGISTERS_reg_24_35_inst : DFF_X1 port map( D => n6316, CK => CLK, Q => 
                           n29479, QN => n18221);
   REGISTERS_reg_24_34_inst : DFF_X1 port map( D => n6315, CK => CLK, Q => 
                           n29478, QN => n18222);
   REGISTERS_reg_24_33_inst : DFF_X1 port map( D => n6314, CK => CLK, Q => 
                           n29477, QN => n18223);
   REGISTERS_reg_24_32_inst : DFF_X1 port map( D => n6313, CK => CLK, Q => 
                           n29476, QN => n18224);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n6312, CK => CLK, Q => 
                           n29475, QN => n18225);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n6311, CK => CLK, Q => 
                           n29474, QN => n18226);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n6310, CK => CLK, Q => 
                           n29473, QN => n18227);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n6309, CK => CLK, Q => 
                           n29472, QN => n18228);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n6308, CK => CLK, Q => 
                           n29471, QN => n18229);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n6307, CK => CLK, Q => 
                           n29470, QN => n18230);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n6306, CK => CLK, Q => 
                           n29469, QN => n18231);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n6305, CK => CLK, Q => 
                           n29468, QN => n18232);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n6304, CK => CLK, Q => 
                           n29467, QN => n18233);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n6303, CK => CLK, Q => 
                           n29466, QN => n18234);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n6302, CK => CLK, Q => 
                           n29465, QN => n18235);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n6301, CK => CLK, Q => 
                           n29464, QN => n18236);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n6300, CK => CLK, Q => 
                           n29463, QN => n18237);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n6299, CK => CLK, Q => 
                           n29462, QN => n18238);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n6298, CK => CLK, Q => 
                           n29461, QN => n18239);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n6297, CK => CLK, Q => 
                           n29460, QN => n18240);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n6296, CK => CLK, Q => 
                           n29459, QN => n18241);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n6295, CK => CLK, Q => 
                           n29458, QN => n18242);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n6294, CK => CLK, Q => 
                           n29457, QN => n18243);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n6293, CK => CLK, Q => 
                           n29456, QN => n18244);
   REGISTERS_reg_14_63_inst : DFF_X1 port map( D => n6984, CK => CLK, Q => 
                           n29635, QN => n17772);
   REGISTERS_reg_14_62_inst : DFF_X1 port map( D => n6983, CK => CLK, Q => 
                           n29634, QN => n17774);
   REGISTERS_reg_14_61_inst : DFF_X1 port map( D => n6982, CK => CLK, Q => 
                           n29633, QN => n17775);
   REGISTERS_reg_14_60_inst : DFF_X1 port map( D => n6981, CK => CLK, Q => 
                           n29632, QN => n17776);
   REGISTERS_reg_14_59_inst : DFF_X1 port map( D => n6980, CK => CLK, Q => 
                           n29631, QN => n17777);
   REGISTERS_reg_14_58_inst : DFF_X1 port map( D => n6979, CK => CLK, Q => 
                           n29630, QN => n17778);
   REGISTERS_reg_14_57_inst : DFF_X1 port map( D => n6978, CK => CLK, Q => 
                           n29629, QN => n17779);
   REGISTERS_reg_14_56_inst : DFF_X1 port map( D => n6977, CK => CLK, Q => 
                           n29628, QN => n17780);
   REGISTERS_reg_14_55_inst : DFF_X1 port map( D => n6976, CK => CLK, Q => 
                           n29627, QN => n17781);
   REGISTERS_reg_14_54_inst : DFF_X1 port map( D => n6975, CK => CLK, Q => 
                           n29626, QN => n17782);
   REGISTERS_reg_14_53_inst : DFF_X1 port map( D => n6974, CK => CLK, Q => 
                           n29625, QN => n17783);
   REGISTERS_reg_14_52_inst : DFF_X1 port map( D => n6973, CK => CLK, Q => 
                           n29624, QN => n17784);
   REGISTERS_reg_14_51_inst : DFF_X1 port map( D => n6972, CK => CLK, Q => 
                           n29623, QN => n17785);
   REGISTERS_reg_14_50_inst : DFF_X1 port map( D => n6971, CK => CLK, Q => 
                           n29622, QN => n17786);
   REGISTERS_reg_14_49_inst : DFF_X1 port map( D => n6970, CK => CLK, Q => 
                           n29621, QN => n17787);
   REGISTERS_reg_14_48_inst : DFF_X1 port map( D => n6969, CK => CLK, Q => 
                           n29620, QN => n17788);
   REGISTERS_reg_14_47_inst : DFF_X1 port map( D => n6968, CK => CLK, Q => 
                           n29619, QN => n17789);
   REGISTERS_reg_14_46_inst : DFF_X1 port map( D => n6967, CK => CLK, Q => 
                           n29618, QN => n17790);
   REGISTERS_reg_14_45_inst : DFF_X1 port map( D => n6966, CK => CLK, Q => 
                           n29617, QN => n17791);
   REGISTERS_reg_14_44_inst : DFF_X1 port map( D => n6965, CK => CLK, Q => 
                           n29616, QN => n17792);
   REGISTERS_reg_14_43_inst : DFF_X1 port map( D => n6964, CK => CLK, Q => 
                           n29615, QN => n17793);
   REGISTERS_reg_14_42_inst : DFF_X1 port map( D => n6963, CK => CLK, Q => 
                           n29614, QN => n17794);
   REGISTERS_reg_14_41_inst : DFF_X1 port map( D => n6962, CK => CLK, Q => 
                           n29613, QN => n17795);
   REGISTERS_reg_14_40_inst : DFF_X1 port map( D => n6961, CK => CLK, Q => 
                           n29612, QN => n17796);
   REGISTERS_reg_14_39_inst : DFF_X1 port map( D => n6960, CK => CLK, Q => 
                           n29611, QN => n17797);
   REGISTERS_reg_14_38_inst : DFF_X1 port map( D => n6959, CK => CLK, Q => 
                           n29610, QN => n17798);
   REGISTERS_reg_14_37_inst : DFF_X1 port map( D => n6958, CK => CLK, Q => 
                           n29609, QN => n17799);
   REGISTERS_reg_14_36_inst : DFF_X1 port map( D => n6957, CK => CLK, Q => 
                           n29608, QN => n17800);
   REGISTERS_reg_14_35_inst : DFF_X1 port map( D => n6956, CK => CLK, Q => 
                           n29607, QN => n17801);
   REGISTERS_reg_14_34_inst : DFF_X1 port map( D => n6955, CK => CLK, Q => 
                           n29606, QN => n17802);
   REGISTERS_reg_14_33_inst : DFF_X1 port map( D => n6954, CK => CLK, Q => 
                           n29605, QN => n17803);
   REGISTERS_reg_14_32_inst : DFF_X1 port map( D => n6953, CK => CLK, Q => 
                           n29604, QN => n17804);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n6952, CK => CLK, Q => 
                           n29603, QN => n17805);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n6951, CK => CLK, Q => 
                           n29602, QN => n17806);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n6950, CK => CLK, Q => 
                           n29601, QN => n17807);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n6949, CK => CLK, Q => 
                           n29600, QN => n17808);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n6948, CK => CLK, Q => 
                           n29599, QN => n17809);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n6947, CK => CLK, Q => 
                           n29598, QN => n17810);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n6946, CK => CLK, Q => 
                           n29597, QN => n17811);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n6945, CK => CLK, Q => 
                           n29596, QN => n17812);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n6944, CK => CLK, Q => 
                           n29595, QN => n17813);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n6943, CK => CLK, Q => 
                           n29594, QN => n17814);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n6942, CK => CLK, Q => 
                           n29593, QN => n17815);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n6941, CK => CLK, Q => 
                           n29592, QN => n17816);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n6940, CK => CLK, Q => 
                           n29591, QN => n17817);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n6939, CK => CLK, Q => 
                           n29590, QN => n17818);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n6938, CK => CLK, Q => 
                           n29589, QN => n17819);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n6937, CK => CLK, Q => 
                           n29588, QN => n17820);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n6936, CK => CLK, Q => 
                           n29587, QN => n17821);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n6935, CK => CLK, Q => 
                           n29586, QN => n17822);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n6934, CK => CLK, Q => 
                           n29585, QN => n17823);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n6933, CK => CLK, Q => 
                           n29584, QN => n17824);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n6932, CK => CLK, Q => 
                           n29583, QN => n17825);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n6931, CK => CLK, Q => 
                           n29582, QN => n17826);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n6930, CK => CLK, Q => 
                           n29581, QN => n17827);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n6929, CK => CLK, Q => 
                           n29580, QN => n17828);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n6928, CK => CLK, Q => 
                           n29579, QN => n17829);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n6927, CK => CLK, Q => 
                           n29578, QN => n17830);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n6926, CK => CLK, Q => 
                           n29577, QN => n17831);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n6925, CK => CLK, Q => 
                           n29576, QN => n17832);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n6924, CK => CLK, Q => 
                           n29575, QN => n17833);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n6923, CK => CLK, Q => 
                           n29574, QN => n17834);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n6922, CK => CLK, Q => 
                           n29573, QN => n17835);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n6921, CK => CLK, Q => 
                           n29572, QN => n17836);
   U13133 : TINV_X1 port map( I => n10761, EN => n5130, ZN => OUT2(63));
   U13134 : TINV_X1 port map( I => n10762, EN => n5132, ZN => OUT2(62));
   U13135 : TINV_X1 port map( I => n10763, EN => n5134, ZN => OUT2(61));
   U13136 : TINV_X1 port map( I => n10764, EN => n5136, ZN => OUT2(60));
   U13137 : TINV_X1 port map( I => n10765, EN => n5138, ZN => OUT2(59));
   U13138 : TINV_X1 port map( I => n10766, EN => n5140, ZN => OUT2(58));
   U13139 : TINV_X1 port map( I => n10767, EN => n5142, ZN => OUT2(57));
   U13140 : TINV_X1 port map( I => n10768, EN => n5144, ZN => OUT2(56));
   U13141 : TINV_X1 port map( I => n10769, EN => n5146, ZN => OUT2(55));
   U13142 : TINV_X1 port map( I => n10770, EN => n5148, ZN => OUT2(54));
   U13143 : TINV_X1 port map( I => n10771, EN => n5150, ZN => OUT2(53));
   U13144 : TINV_X1 port map( I => n10772, EN => n5152, ZN => OUT2(52));
   U13145 : TINV_X1 port map( I => n10773, EN => n5154, ZN => OUT2(51));
   U13146 : TINV_X1 port map( I => n10774, EN => n5156, ZN => OUT2(50));
   U13147 : TINV_X1 port map( I => n10775, EN => n5158, ZN => OUT2(49));
   U13148 : TINV_X1 port map( I => n10776, EN => n5160, ZN => OUT2(48));
   U13149 : TINV_X1 port map( I => n10777, EN => n5162, ZN => OUT2(47));
   U13150 : TINV_X1 port map( I => n10778, EN => n5164, ZN => OUT2(46));
   U13151 : TINV_X1 port map( I => n10779, EN => n5166, ZN => OUT2(45));
   U13152 : TINV_X1 port map( I => n10780, EN => n5168, ZN => OUT2(44));
   U13153 : TINV_X1 port map( I => n10781, EN => n5170, ZN => OUT2(43));
   U13154 : TINV_X1 port map( I => n10782, EN => n5172, ZN => OUT2(42));
   U13155 : TINV_X1 port map( I => n10783, EN => n5174, ZN => OUT2(41));
   U13156 : TINV_X1 port map( I => n10784, EN => n5176, ZN => OUT2(40));
   U13157 : TINV_X1 port map( I => n10785, EN => n5178, ZN => OUT2(39));
   U13158 : TINV_X1 port map( I => n10786, EN => n5180, ZN => OUT2(38));
   U13159 : TINV_X1 port map( I => n10787, EN => n5182, ZN => OUT2(37));
   U13160 : TINV_X1 port map( I => n10788, EN => n5184, ZN => OUT2(36));
   U13161 : TINV_X1 port map( I => n10789, EN => n5186, ZN => OUT2(35));
   U13162 : TINV_X1 port map( I => n10790, EN => n5188, ZN => OUT2(34));
   U13163 : TINV_X1 port map( I => n10791, EN => n5190, ZN => OUT2(33));
   U13164 : TINV_X1 port map( I => n10792, EN => n5192, ZN => OUT2(32));
   U13165 : TINV_X1 port map( I => n10793, EN => n5194, ZN => OUT2(31));
   U13166 : TINV_X1 port map( I => n10794, EN => n5196, ZN => OUT2(30));
   U13167 : TINV_X1 port map( I => n10795, EN => n5198, ZN => OUT2(29));
   U13168 : TINV_X1 port map( I => n10796, EN => n5200, ZN => OUT2(28));
   U13169 : TINV_X1 port map( I => n10797, EN => n5202, ZN => OUT2(27));
   U13170 : TINV_X1 port map( I => n10798, EN => n5204, ZN => OUT2(26));
   U13171 : TINV_X1 port map( I => n10799, EN => n5206, ZN => OUT2(25));
   U13172 : TINV_X1 port map( I => n10800, EN => n5208, ZN => OUT2(24));
   U13173 : TINV_X1 port map( I => n10801, EN => n5210, ZN => OUT2(23));
   U13174 : TINV_X1 port map( I => n10802, EN => n5212, ZN => OUT2(22));
   U13175 : TINV_X1 port map( I => n10803, EN => n5214, ZN => OUT2(21));
   U13176 : TINV_X1 port map( I => n10804, EN => n5216, ZN => OUT2(20));
   U13177 : TINV_X1 port map( I => n10805, EN => n5218, ZN => OUT2(19));
   U13178 : TINV_X1 port map( I => n10806, EN => n5220, ZN => OUT2(18));
   U13179 : TINV_X1 port map( I => n10807, EN => n5222, ZN => OUT2(17));
   U13180 : TINV_X1 port map( I => n10808, EN => n5224, ZN => OUT2(16));
   U13181 : TINV_X1 port map( I => n10809, EN => n5226, ZN => OUT2(15));
   U13182 : TINV_X1 port map( I => n10810, EN => n5228, ZN => OUT2(14));
   U13183 : TINV_X1 port map( I => n10811, EN => n5230, ZN => OUT2(13));
   U13184 : TINV_X1 port map( I => n10812, EN => n5232, ZN => OUT2(12));
   U13185 : TINV_X1 port map( I => n10813, EN => n5234, ZN => OUT2(11));
   U13186 : TINV_X1 port map( I => n10814, EN => n5236, ZN => OUT2(10));
   U13187 : TINV_X1 port map( I => n10815, EN => n5238, ZN => OUT2(9));
   U13188 : TINV_X1 port map( I => n10816, EN => n5240, ZN => OUT2(8));
   U13189 : TINV_X1 port map( I => n10817, EN => n5242, ZN => OUT2(7));
   U13190 : TINV_X1 port map( I => n10818, EN => n5244, ZN => OUT2(6));
   U13191 : TINV_X1 port map( I => n10819, EN => n5246, ZN => OUT2(5));
   U13192 : TINV_X1 port map( I => n10820, EN => n5248, ZN => OUT2(4));
   U13193 : TINV_X1 port map( I => n10821, EN => n5250, ZN => OUT2(3));
   U13194 : TINV_X1 port map( I => n10822, EN => n5252, ZN => OUT2(2));
   U13195 : TINV_X1 port map( I => n10823, EN => n5254, ZN => OUT2(1));
   U13196 : TINV_X1 port map( I => n10824, EN => n5256, ZN => OUT2(0));
   U13197 : TINV_X1 port map( I => n10825, EN => n5258, ZN => OUT1(63));
   U13198 : TINV_X1 port map( I => n10826, EN => n5260, ZN => OUT1(62));
   U13199 : TINV_X1 port map( I => n10827, EN => n5262, ZN => OUT1(61));
   U13200 : TINV_X1 port map( I => n10828, EN => n5264, ZN => OUT1(60));
   U13201 : TINV_X1 port map( I => n10829, EN => n5266, ZN => OUT1(59));
   U13202 : TINV_X1 port map( I => n10830, EN => n5268, ZN => OUT1(58));
   U13203 : TINV_X1 port map( I => n10831, EN => n5270, ZN => OUT1(57));
   U13204 : TINV_X1 port map( I => n10832, EN => n5272, ZN => OUT1(56));
   U13205 : TINV_X1 port map( I => n10833, EN => n5274, ZN => OUT1(55));
   U13206 : TINV_X1 port map( I => n10834, EN => n5276, ZN => OUT1(54));
   U13207 : TINV_X1 port map( I => n10835, EN => n5278, ZN => OUT1(53));
   U13208 : TINV_X1 port map( I => n10836, EN => n5280, ZN => OUT1(52));
   U13209 : TINV_X1 port map( I => n10837, EN => n5282, ZN => OUT1(51));
   U13210 : TINV_X1 port map( I => n10838, EN => n5284, ZN => OUT1(50));
   U13211 : TINV_X1 port map( I => n10839, EN => n5286, ZN => OUT1(49));
   U13212 : TINV_X1 port map( I => n10840, EN => n5288, ZN => OUT1(48));
   U13213 : TINV_X1 port map( I => n10841, EN => n5290, ZN => OUT1(47));
   U13214 : TINV_X1 port map( I => n10842, EN => n5292, ZN => OUT1(46));
   U13215 : TINV_X1 port map( I => n10843, EN => n5294, ZN => OUT1(45));
   U13216 : TINV_X1 port map( I => n10844, EN => n5296, ZN => OUT1(44));
   U13217 : TINV_X1 port map( I => n10845, EN => n5298, ZN => OUT1(43));
   U13218 : TINV_X1 port map( I => n10846, EN => n5300, ZN => OUT1(42));
   U13219 : TINV_X1 port map( I => n10847, EN => n5302, ZN => OUT1(41));
   U13220 : TINV_X1 port map( I => n10848, EN => n5304, ZN => OUT1(40));
   U13221 : TINV_X1 port map( I => n10849, EN => n5306, ZN => OUT1(39));
   U13222 : TINV_X1 port map( I => n10850, EN => n5308, ZN => OUT1(38));
   U13223 : TINV_X1 port map( I => n10851, EN => n5310, ZN => OUT1(37));
   U13224 : TINV_X1 port map( I => n10852, EN => n5312, ZN => OUT1(36));
   U13225 : TINV_X1 port map( I => n10853, EN => n5314, ZN => OUT1(35));
   U13226 : TINV_X1 port map( I => n10854, EN => n5316, ZN => OUT1(34));
   U13227 : TINV_X1 port map( I => n10855, EN => n5318, ZN => OUT1(33));
   U13228 : TINV_X1 port map( I => n10856, EN => n5320, ZN => OUT1(32));
   U13229 : TINV_X1 port map( I => n10857, EN => n5322, ZN => OUT1(31));
   U13230 : TINV_X1 port map( I => n10858, EN => n5324, ZN => OUT1(30));
   U13231 : TINV_X1 port map( I => n10859, EN => n5326, ZN => OUT1(29));
   U13232 : TINV_X1 port map( I => n10860, EN => n5328, ZN => OUT1(28));
   U13233 : TINV_X1 port map( I => n10861, EN => n5330, ZN => OUT1(27));
   U13234 : TINV_X1 port map( I => n10862, EN => n5332, ZN => OUT1(26));
   U13235 : TINV_X1 port map( I => n10863, EN => n5334, ZN => OUT1(25));
   U13236 : TINV_X1 port map( I => n10864, EN => n5336, ZN => OUT1(24));
   U13237 : TINV_X1 port map( I => n10865, EN => n5338, ZN => OUT1(23));
   U13238 : TINV_X1 port map( I => n10866, EN => n5340, ZN => OUT1(22));
   U13239 : TINV_X1 port map( I => n10867, EN => n5342, ZN => OUT1(21));
   U13240 : TINV_X1 port map( I => n10868, EN => n5344, ZN => OUT1(20));
   U13241 : TINV_X1 port map( I => n10869, EN => n5346, ZN => OUT1(19));
   U13242 : TINV_X1 port map( I => n10870, EN => n5348, ZN => OUT1(18));
   U13243 : TINV_X1 port map( I => n10871, EN => n5350, ZN => OUT1(17));
   U13244 : TINV_X1 port map( I => n10872, EN => n5352, ZN => OUT1(16));
   U13245 : TINV_X1 port map( I => n10873, EN => n5354, ZN => OUT1(15));
   U13246 : TINV_X1 port map( I => n10874, EN => n5356, ZN => OUT1(14));
   U13247 : TINV_X1 port map( I => n10875, EN => n5358, ZN => OUT1(13));
   U13248 : TINV_X1 port map( I => n10876, EN => n5360, ZN => OUT1(12));
   U13249 : TINV_X1 port map( I => n10877, EN => n5362, ZN => OUT1(11));
   U13250 : TINV_X1 port map( I => n10878, EN => n5364, ZN => OUT1(10));
   U13251 : TINV_X1 port map( I => n10879, EN => n5366, ZN => OUT1(9));
   U13252 : TINV_X1 port map( I => n10880, EN => n5368, ZN => OUT1(8));
   U13253 : TINV_X1 port map( I => n10881, EN => n5370, ZN => OUT1(7));
   U13254 : TINV_X1 port map( I => n10882, EN => n5372, ZN => OUT1(6));
   U13255 : TINV_X1 port map( I => n10883, EN => n5374, ZN => OUT1(5));
   U13256 : TINV_X1 port map( I => n10884, EN => n5376, ZN => OUT1(4));
   U13257 : TINV_X1 port map( I => n10885, EN => n5378, ZN => OUT1(3));
   U13258 : TINV_X1 port map( I => n10886, EN => n5380, ZN => OUT1(2));
   U13259 : TINV_X1 port map( I => n10887, EN => n5382, ZN => OUT1(1));
   U13260 : TINV_X1 port map( I => n10888, EN => n5384, ZN => OUT1(0));
   U19722 : NAND3_X1 port map( A1 => n25452, A2 => n25453, A3 => n25454, ZN => 
                           n25231);
   U19723 : NAND3_X1 port map( A1 => n25454, A2 => n25453, A3 => ADD_WR(0), ZN 
                           => n25235);
   U19724 : NAND3_X1 port map( A1 => n25454, A2 => n25452, A3 => ADD_WR(3), ZN 
                           => n25587);
   U19725 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n25454, A3 => ADD_WR(3), 
                           ZN => n25654);
   U19726 : NAND3_X1 port map( A1 => n25452, A2 => n25453, A3 => n26091, ZN => 
                           n25873);
   U19727 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n25453, A3 => n26091, ZN 
                           => n25940);
   U19728 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => n25452, A3 => n26091, ZN 
                           => n26096);
   U19729 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => ADD_WR(0), A3 => n26091, 
                           ZN => n26099);
   REGISTERS_reg_30_63_inst : DFF_X1 port map( D => n5960, CK => CLK, Q => 
                           n30140, QN => n26251);
   REGISTERS_reg_30_62_inst : DFF_X1 port map( D => n5959, CK => CLK, Q => 
                           n30139, QN => n26253);
   REGISTERS_reg_30_61_inst : DFF_X1 port map( D => n5958, CK => CLK, Q => 
                           n30138, QN => n26254);
   REGISTERS_reg_30_60_inst : DFF_X1 port map( D => n5957, CK => CLK, Q => 
                           n30137, QN => n26255);
   REGISTERS_reg_27_63_inst : DFF_X1 port map( D => n6152, CK => CLK, Q => 
                           n22011, QN => n26169);
   REGISTERS_reg_27_62_inst : DFF_X1 port map( D => n6151, CK => CLK, Q => 
                           n22010, QN => n26171);
   REGISTERS_reg_27_61_inst : DFF_X1 port map( D => n6150, CK => CLK, Q => 
                           n22009, QN => n26172);
   REGISTERS_reg_27_60_inst : DFF_X1 port map( D => n6149, CK => CLK, Q => 
                           n22008, QN => n26173);
   REGISTERS_reg_26_63_inst : DFF_X1 port map( D => n6216, CK => CLK, Q => 
                           n9292, QN => n26103);
   REGISTERS_reg_26_62_inst : DFF_X1 port map( D => n6215, CK => CLK, Q => 
                           n9297, QN => n26105);
   REGISTERS_reg_26_61_inst : DFF_X1 port map( D => n6214, CK => CLK, Q => 
                           n9302, QN => n26106);
   REGISTERS_reg_26_60_inst : DFF_X1 port map( D => n6213, CK => CLK, Q => 
                           n9307, QN => n26107);
   REGISTERS_reg_21_63_inst : DFF_X1 port map( D => n6536, CK => CLK, Q => 
                           n30136, QN => n26024);
   REGISTERS_reg_21_62_inst : DFF_X1 port map( D => n6535, CK => CLK, Q => 
                           n30135, QN => n26026);
   REGISTERS_reg_21_61_inst : DFF_X1 port map( D => n6534, CK => CLK, Q => 
                           n30134, QN => n26027);
   REGISTERS_reg_21_60_inst : DFF_X1 port map( D => n6533, CK => CLK, Q => 
                           n30133, QN => n26028);
   REGISTERS_reg_20_63_inst : DFF_X1 port map( D => n6600, CK => CLK, Q => 
                           n30132, QN => n25958);
   REGISTERS_reg_20_62_inst : DFF_X1 port map( D => n6599, CK => CLK, Q => 
                           n30131, QN => n25960);
   REGISTERS_reg_20_61_inst : DFF_X1 port map( D => n6598, CK => CLK, Q => 
                           n30130, QN => n25961);
   REGISTERS_reg_20_60_inst : DFF_X1 port map( D => n6597, CK => CLK, Q => 
                           n30129, QN => n25962);
   REGISTERS_reg_16_63_inst : DFF_X1 port map( D => n6856, CK => CLK, Q => 
                           n9293, QN => n25808);
   REGISTERS_reg_16_62_inst : DFF_X1 port map( D => n6855, CK => CLK, Q => 
                           n9298, QN => n25810);
   REGISTERS_reg_16_61_inst : DFF_X1 port map( D => n6854, CK => CLK, Q => 
                           n9303, QN => n25811);
   REGISTERS_reg_16_60_inst : DFF_X1 port map( D => n6853, CK => CLK, Q => 
                           n9308, QN => n25812);
   REGISTERS_reg_17_63_inst : DFF_X1 port map( D => n6792, CK => CLK, Q => 
                           n21922, QN => n25875);
   REGISTERS_reg_17_62_inst : DFF_X1 port map( D => n6791, CK => CLK, Q => 
                           n21921, QN => n25877);
   REGISTERS_reg_17_61_inst : DFF_X1 port map( D => n6790, CK => CLK, Q => 
                           n21920, QN => n25878);
   REGISTERS_reg_17_60_inst : DFF_X1 port map( D => n6789, CK => CLK, Q => 
                           n21919, QN => n25879);
   REGISTERS_reg_31_63_inst : DFF_X1 port map( D => n5896, CK => CLK, Q => 
                           n30128, QN => n26317);
   REGISTERS_reg_31_62_inst : DFF_X1 port map( D => n5894, CK => CLK, Q => 
                           n30127, QN => n26378);
   REGISTERS_reg_31_61_inst : DFF_X1 port map( D => n5892, CK => CLK, Q => 
                           n30126, QN => n26404);
   REGISTERS_reg_31_60_inst : DFF_X1 port map( D => n5890, CK => CLK, Q => 
                           n30125, QN => n26430);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n6028, CK => CLK, Q => 
                           n30124, QN => n26244);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n6027, CK => CLK, Q => 
                           n30123, QN => n26245);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n6026, CK => CLK, Q => 
                           n30122, QN => n26246);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n6025, CK => CLK, Q => 
                           n30121, QN => n26247);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n6668, CK => CLK, Q => 
                           n30120, QN => n25951);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n6667, CK => CLK, Q => 
                           n30119, QN => n25952);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n6666, CK => CLK, Q => 
                           n30118, QN => n25953);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n6665, CK => CLK, Q => 
                           n30117, QN => n25954);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n6036, CK => CLK, Q => 
                           n30116, QN => n26236);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n6035, CK => CLK, Q => 
                           n30115, QN => n26237);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n6034, CK => CLK, Q => 
                           n30114, QN => n26238);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n6033, CK => CLK, Q => 
                           n30113, QN => n26239);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n6032, CK => CLK, Q => 
                           n30112, QN => n26240);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n6031, CK => CLK, Q => 
                           n30111, QN => n26241);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n6030, CK => CLK, Q => 
                           n30110, QN => n26242);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n6029, CK => CLK, Q => 
                           n30109, QN => n26243);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n6676, CK => CLK, Q => 
                           n30108, QN => n25943);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n6675, CK => CLK, Q => 
                           n30107, QN => n25944);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n6674, CK => CLK, Q => 
                           n30106, QN => n25945);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n6673, CK => CLK, Q => 
                           n30105, QN => n25946);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n6672, CK => CLK, Q => 
                           n30104, QN => n25947);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n6671, CK => CLK, Q => 
                           n30103, QN => n25948);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n6670, CK => CLK, Q => 
                           n30102, QN => n25949);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n6669, CK => CLK, Q => 
                           n30101, QN => n25950);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n5792, CK => CLK, Q => 
                           n30100, QN => n27704);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n5790, CK => CLK, Q => 
                           n30099, QN => n27730);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n5788, CK => CLK, Q => 
                           n30098, QN => n27756);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n5786, CK => CLK, Q => 
                           n30097, QN => n27782);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n5784, CK => CLK, Q => 
                           n30096, QN => n27808);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n5782, CK => CLK, Q => 
                           n30095, QN => n27834);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n5780, CK => CLK, Q => 
                           n30094, QN => n27860);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n5778, CK => CLK, Q => 
                           n30093, QN => n27886);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n5776, CK => CLK, Q => 
                           n30092, QN => n27912);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n5774, CK => CLK, Q => 
                           n30091, QN => n27938);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n5772, CK => CLK, Q => 
                           n30090, QN => n27964);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n5770, CK => CLK, Q => 
                           n30089, QN => n27990);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n5908, CK => CLK, Q => 
                           n30088, QN => n26304);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n5907, CK => CLK, Q => 
                           n30087, QN => n26305);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n5906, CK => CLK, Q => 
                           n30086, QN => n26306);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n5905, CK => CLK, Q => 
                           n30085, QN => n26307);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n5904, CK => CLK, Q => 
                           n30084, QN => n26308);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n5903, CK => CLK, Q => 
                           n30083, QN => n26309);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n5902, CK => CLK, Q => 
                           n30082, QN => n26310);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n5901, CK => CLK, Q => 
                           n30081, QN => n26311);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n5900, CK => CLK, Q => 
                           n30080, QN => n26312);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n5899, CK => CLK, Q => 
                           n30079, QN => n26313);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n5898, CK => CLK, Q => 
                           n30078, QN => n26314);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n5897, CK => CLK, Q => 
                           n30077, QN => n26315);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n6100, CK => CLK, Q => 
                           n21998, QN => n26222);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n6099, CK => CLK, Q => 
                           n21997, QN => n26223);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n6098, CK => CLK, Q => 
                           n21996, QN => n26224);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n6097, CK => CLK, Q => 
                           n21995, QN => n26225);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n6096, CK => CLK, Q => 
                           n21994, QN => n26226);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n6095, CK => CLK, Q => 
                           n21993, QN => n26227);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n6094, CK => CLK, Q => 
                           n21992, QN => n26228);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n6093, CK => CLK, Q => 
                           n21991, QN => n26229);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n6092, CK => CLK, Q => 
                           n21990, QN => n26230);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n6091, CK => CLK, Q => 
                           n21989, QN => n26231);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n6090, CK => CLK, Q => 
                           n21988, QN => n26232);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n6089, CK => CLK, Q => 
                           n21987, QN => n26233);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n6164, CK => CLK, Q => 
                           n9552, QN => n26156);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n6163, CK => CLK, Q => 
                           n9557, QN => n26157);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n6162, CK => CLK, Q => n9562
                           , QN => n26158);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n6161, CK => CLK, Q => n9567
                           , QN => n26159);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n6160, CK => CLK, Q => n9572
                           , QN => n26160);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n6159, CK => CLK, Q => n9577
                           , QN => n26161);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n6158, CK => CLK, Q => n9582
                           , QN => n26162);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n6157, CK => CLK, Q => n9587
                           , QN => n26163);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n6156, CK => CLK, Q => n9592
                           , QN => n26164);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n6155, CK => CLK, Q => n9597
                           , QN => n26165);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n6154, CK => CLK, Q => n9602
                           , QN => n26166);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n6153, CK => CLK, Q => n9607
                           , QN => n26167);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n6484, CK => CLK, Q => 
                           n30076, QN => n26077);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n6483, CK => CLK, Q => 
                           n30075, QN => n26078);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n6482, CK => CLK, Q => 
                           n30074, QN => n26079);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n6481, CK => CLK, Q => 
                           n30073, QN => n26080);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n6480, CK => CLK, Q => 
                           n30072, QN => n26081);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n6479, CK => CLK, Q => 
                           n30071, QN => n26082);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n6478, CK => CLK, Q => 
                           n30070, QN => n26083);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n6477, CK => CLK, Q => 
                           n30069, QN => n26084);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n6476, CK => CLK, Q => 
                           n30068, QN => n26085);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n6475, CK => CLK, Q => 
                           n30067, QN => n26086);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n6474, CK => CLK, Q => 
                           n30066, QN => n26087);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n6473, CK => CLK, Q => 
                           n30065, QN => n26088);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n6548, CK => CLK, Q => 
                           n30064, QN => n26011);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n6547, CK => CLK, Q => 
                           n30063, QN => n26012);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n6546, CK => CLK, Q => 
                           n30062, QN => n26013);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n6545, CK => CLK, Q => 
                           n30061, QN => n26014);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n6544, CK => CLK, Q => 
                           n30060, QN => n26015);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n6543, CK => CLK, Q => 
                           n30059, QN => n26016);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n6542, CK => CLK, Q => 
                           n30058, QN => n26017);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n6541, CK => CLK, Q => 
                           n30057, QN => n26018);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n6540, CK => CLK, Q => 
                           n30056, QN => n26019);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n6539, CK => CLK, Q => 
                           n30055, QN => n26020);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n6538, CK => CLK, Q => 
                           n30054, QN => n26021);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n6537, CK => CLK, Q => 
                           n30053, QN => n26022);
   REGISTERS_reg_31_59_inst : DFF_X1 port map( D => n5888, CK => CLK, Q => 
                           n30052, QN => n26456);
   REGISTERS_reg_31_58_inst : DFF_X1 port map( D => n5886, CK => CLK, Q => 
                           n30051, QN => n26482);
   REGISTERS_reg_31_57_inst : DFF_X1 port map( D => n5884, CK => CLK, Q => 
                           n30050, QN => n26508);
   REGISTERS_reg_31_56_inst : DFF_X1 port map( D => n5882, CK => CLK, Q => 
                           n30049, QN => n26534);
   REGISTERS_reg_31_55_inst : DFF_X1 port map( D => n5880, CK => CLK, Q => 
                           n30048, QN => n26560);
   REGISTERS_reg_31_54_inst : DFF_X1 port map( D => n5878, CK => CLK, Q => 
                           n30047, QN => n26586);
   REGISTERS_reg_31_53_inst : DFF_X1 port map( D => n5876, CK => CLK, Q => 
                           n30046, QN => n26612);
   REGISTERS_reg_31_52_inst : DFF_X1 port map( D => n5874, CK => CLK, Q => 
                           n30045, QN => n26638);
   REGISTERS_reg_31_51_inst : DFF_X1 port map( D => n5872, CK => CLK, Q => 
                           n30044, QN => n26664);
   REGISTERS_reg_31_50_inst : DFF_X1 port map( D => n5870, CK => CLK, Q => 
                           n30043, QN => n26690);
   REGISTERS_reg_31_49_inst : DFF_X1 port map( D => n5868, CK => CLK, Q => 
                           n30042, QN => n26716);
   REGISTERS_reg_31_48_inst : DFF_X1 port map( D => n5866, CK => CLK, Q => 
                           n30041, QN => n26742);
   REGISTERS_reg_31_47_inst : DFF_X1 port map( D => n5864, CK => CLK, Q => 
                           n30040, QN => n26768);
   REGISTERS_reg_31_46_inst : DFF_X1 port map( D => n5862, CK => CLK, Q => 
                           n30039, QN => n26794);
   REGISTERS_reg_31_45_inst : DFF_X1 port map( D => n5860, CK => CLK, Q => 
                           n30038, QN => n26820);
   REGISTERS_reg_31_44_inst : DFF_X1 port map( D => n5858, CK => CLK, Q => 
                           n30037, QN => n26846);
   REGISTERS_reg_31_43_inst : DFF_X1 port map( D => n5856, CK => CLK, Q => 
                           n30036, QN => n26872);
   REGISTERS_reg_31_42_inst : DFF_X1 port map( D => n5854, CK => CLK, Q => 
                           n30035, QN => n26898);
   REGISTERS_reg_31_41_inst : DFF_X1 port map( D => n5852, CK => CLK, Q => 
                           n30034, QN => n26924);
   REGISTERS_reg_31_40_inst : DFF_X1 port map( D => n5850, CK => CLK, Q => 
                           n30033, QN => n26950);
   REGISTERS_reg_31_39_inst : DFF_X1 port map( D => n5848, CK => CLK, Q => 
                           n30032, QN => n26976);
   REGISTERS_reg_31_38_inst : DFF_X1 port map( D => n5846, CK => CLK, Q => 
                           n30031, QN => n27002);
   REGISTERS_reg_31_37_inst : DFF_X1 port map( D => n5844, CK => CLK, Q => 
                           n30030, QN => n27028);
   REGISTERS_reg_31_36_inst : DFF_X1 port map( D => n5842, CK => CLK, Q => 
                           n30029, QN => n27054);
   REGISTERS_reg_31_35_inst : DFF_X1 port map( D => n5840, CK => CLK, Q => 
                           n30028, QN => n27080);
   REGISTERS_reg_31_34_inst : DFF_X1 port map( D => n5838, CK => CLK, Q => 
                           n30027, QN => n27106);
   REGISTERS_reg_31_33_inst : DFF_X1 port map( D => n5836, CK => CLK, Q => 
                           n30026, QN => n27132);
   REGISTERS_reg_31_32_inst : DFF_X1 port map( D => n5834, CK => CLK, Q => 
                           n30025, QN => n27158);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n5832, CK => CLK, Q => 
                           n30024, QN => n27184);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n5830, CK => CLK, Q => 
                           n30023, QN => n27210);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n5828, CK => CLK, Q => 
                           n30022, QN => n27236);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n5826, CK => CLK, Q => 
                           n30021, QN => n27262);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n5824, CK => CLK, Q => 
                           n30020, QN => n27288);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n5822, CK => CLK, Q => 
                           n30019, QN => n27314);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n5820, CK => CLK, Q => 
                           n30018, QN => n27340);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n5818, CK => CLK, Q => 
                           n30017, QN => n27366);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n5816, CK => CLK, Q => 
                           n30016, QN => n27392);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n5814, CK => CLK, Q => 
                           n30015, QN => n27418);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n5812, CK => CLK, Q => 
                           n30014, QN => n27444);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n5810, CK => CLK, Q => 
                           n30013, QN => n27470);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n5808, CK => CLK, Q => 
                           n30012, QN => n27496);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n5806, CK => CLK, Q => 
                           n30011, QN => n27522);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n5804, CK => CLK, Q => 
                           n30010, QN => n27548);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n5802, CK => CLK, Q => 
                           n30009, QN => n27574);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n5800, CK => CLK, Q => 
                           n30008, QN => n27600);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n5798, CK => CLK, Q => 
                           n30007, QN => n27626);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n5796, CK => CLK, Q => 
                           n30006, QN => n27652);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n5794, CK => CLK, Q => 
                           n30005, QN => n27678);
   REGISTERS_reg_30_59_inst : DFF_X1 port map( D => n5956, CK => CLK, Q => 
                           n30004, QN => n26256);
   REGISTERS_reg_30_58_inst : DFF_X1 port map( D => n5955, CK => CLK, Q => 
                           n30003, QN => n26257);
   REGISTERS_reg_30_57_inst : DFF_X1 port map( D => n5954, CK => CLK, Q => 
                           n30002, QN => n26258);
   REGISTERS_reg_30_56_inst : DFF_X1 port map( D => n5953, CK => CLK, Q => 
                           n30001, QN => n26259);
   REGISTERS_reg_30_55_inst : DFF_X1 port map( D => n5952, CK => CLK, Q => 
                           n30000, QN => n26260);
   REGISTERS_reg_30_54_inst : DFF_X1 port map( D => n5951, CK => CLK, Q => 
                           n29999, QN => n26261);
   REGISTERS_reg_30_53_inst : DFF_X1 port map( D => n5950, CK => CLK, Q => 
                           n29998, QN => n26262);
   REGISTERS_reg_30_52_inst : DFF_X1 port map( D => n5949, CK => CLK, Q => 
                           n29997, QN => n26263);
   REGISTERS_reg_30_51_inst : DFF_X1 port map( D => n5948, CK => CLK, Q => 
                           n29996, QN => n26264);
   REGISTERS_reg_30_50_inst : DFF_X1 port map( D => n5947, CK => CLK, Q => 
                           n29995, QN => n26265);
   REGISTERS_reg_30_49_inst : DFF_X1 port map( D => n5946, CK => CLK, Q => 
                           n29994, QN => n26266);
   REGISTERS_reg_30_48_inst : DFF_X1 port map( D => n5945, CK => CLK, Q => 
                           n29993, QN => n26267);
   REGISTERS_reg_30_47_inst : DFF_X1 port map( D => n5944, CK => CLK, Q => 
                           n29992, QN => n26268);
   REGISTERS_reg_30_46_inst : DFF_X1 port map( D => n5943, CK => CLK, Q => 
                           n29991, QN => n26269);
   REGISTERS_reg_30_45_inst : DFF_X1 port map( D => n5942, CK => CLK, Q => 
                           n29990, QN => n26270);
   REGISTERS_reg_30_44_inst : DFF_X1 port map( D => n5941, CK => CLK, Q => 
                           n29989, QN => n26271);
   REGISTERS_reg_30_43_inst : DFF_X1 port map( D => n5940, CK => CLK, Q => 
                           n29988, QN => n26272);
   REGISTERS_reg_30_42_inst : DFF_X1 port map( D => n5939, CK => CLK, Q => 
                           n29987, QN => n26273);
   REGISTERS_reg_30_41_inst : DFF_X1 port map( D => n5938, CK => CLK, Q => 
                           n29986, QN => n26274);
   REGISTERS_reg_30_40_inst : DFF_X1 port map( D => n5937, CK => CLK, Q => 
                           n29985, QN => n26275);
   REGISTERS_reg_30_39_inst : DFF_X1 port map( D => n5936, CK => CLK, Q => 
                           n29984, QN => n26276);
   REGISTERS_reg_30_38_inst : DFF_X1 port map( D => n5935, CK => CLK, Q => 
                           n29983, QN => n26277);
   REGISTERS_reg_30_37_inst : DFF_X1 port map( D => n5934, CK => CLK, Q => 
                           n29982, QN => n26278);
   REGISTERS_reg_30_36_inst : DFF_X1 port map( D => n5933, CK => CLK, Q => 
                           n29981, QN => n26279);
   REGISTERS_reg_30_35_inst : DFF_X1 port map( D => n5932, CK => CLK, Q => 
                           n29980, QN => n26280);
   REGISTERS_reg_30_34_inst : DFF_X1 port map( D => n5931, CK => CLK, Q => 
                           n29979, QN => n26281);
   REGISTERS_reg_30_33_inst : DFF_X1 port map( D => n5930, CK => CLK, Q => 
                           n29978, QN => n26282);
   REGISTERS_reg_30_32_inst : DFF_X1 port map( D => n5929, CK => CLK, Q => 
                           n29977, QN => n26283);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n5928, CK => CLK, Q => 
                           n29976, QN => n26284);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n5927, CK => CLK, Q => 
                           n29975, QN => n26285);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n5926, CK => CLK, Q => 
                           n29974, QN => n26286);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n5925, CK => CLK, Q => 
                           n29973, QN => n26287);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n5924, CK => CLK, Q => 
                           n29972, QN => n26288);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n5923, CK => CLK, Q => 
                           n29971, QN => n26289);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n5922, CK => CLK, Q => 
                           n29970, QN => n26290);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n5921, CK => CLK, Q => 
                           n29969, QN => n26291);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n5920, CK => CLK, Q => 
                           n29968, QN => n26292);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n5919, CK => CLK, Q => 
                           n29967, QN => n26293);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n5918, CK => CLK, Q => 
                           n29966, QN => n26294);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n5917, CK => CLK, Q => 
                           n29965, QN => n26295);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n5916, CK => CLK, Q => 
                           n29964, QN => n26296);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n5915, CK => CLK, Q => 
                           n29963, QN => n26297);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n5914, CK => CLK, Q => 
                           n29962, QN => n26298);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n5913, CK => CLK, Q => 
                           n29961, QN => n26299);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n5912, CK => CLK, Q => 
                           n29960, QN => n26300);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n5911, CK => CLK, Q => 
                           n29959, QN => n26301);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n5910, CK => CLK, Q => 
                           n29958, QN => n26302);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n5909, CK => CLK, Q => 
                           n29957, QN => n26303);
   REGISTERS_reg_27_59_inst : DFF_X1 port map( D => n6148, CK => CLK, Q => 
                           n22007, QN => n26174);
   REGISTERS_reg_27_58_inst : DFF_X1 port map( D => n6147, CK => CLK, Q => 
                           n22006, QN => n26175);
   REGISTERS_reg_27_57_inst : DFF_X1 port map( D => n6146, CK => CLK, Q => 
                           n22005, QN => n26176);
   REGISTERS_reg_27_56_inst : DFF_X1 port map( D => n6145, CK => CLK, Q => 
                           n22004, QN => n26177);
   REGISTERS_reg_27_55_inst : DFF_X1 port map( D => n6144, CK => CLK, Q => 
                           n22003, QN => n26178);
   REGISTERS_reg_27_54_inst : DFF_X1 port map( D => n6143, CK => CLK, Q => 
                           n22002, QN => n26179);
   REGISTERS_reg_27_53_inst : DFF_X1 port map( D => n6142, CK => CLK, Q => 
                           n22001, QN => n26180);
   REGISTERS_reg_27_52_inst : DFF_X1 port map( D => n6141, CK => CLK, Q => 
                           n22000, QN => n26181);
   REGISTERS_reg_27_51_inst : DFF_X1 port map( D => n6140, CK => CLK, Q => 
                           n21999, QN => n26182);
   REGISTERS_reg_27_50_inst : DFF_X1 port map( D => n6139, CK => CLK, Q => 
                           n22114, QN => n26183);
   REGISTERS_reg_27_49_inst : DFF_X1 port map( D => n6138, CK => CLK, Q => 
                           n22113, QN => n26184);
   REGISTERS_reg_27_48_inst : DFF_X1 port map( D => n6137, CK => CLK, Q => 
                           n22112, QN => n26185);
   REGISTERS_reg_27_47_inst : DFF_X1 port map( D => n6136, CK => CLK, Q => 
                           n22111, QN => n26186);
   REGISTERS_reg_27_46_inst : DFF_X1 port map( D => n6135, CK => CLK, Q => 
                           n22110, QN => n26187);
   REGISTERS_reg_27_45_inst : DFF_X1 port map( D => n6134, CK => CLK, Q => 
                           n22109, QN => n26188);
   REGISTERS_reg_27_44_inst : DFF_X1 port map( D => n6133, CK => CLK, Q => 
                           n22108, QN => n26189);
   REGISTERS_reg_27_43_inst : DFF_X1 port map( D => n6132, CK => CLK, Q => 
                           n22107, QN => n26190);
   REGISTERS_reg_27_42_inst : DFF_X1 port map( D => n6131, CK => CLK, Q => 
                           n22106, QN => n26191);
   REGISTERS_reg_27_41_inst : DFF_X1 port map( D => n6130, CK => CLK, Q => 
                           n22105, QN => n26192);
   REGISTERS_reg_27_40_inst : DFF_X1 port map( D => n6129, CK => CLK, Q => 
                           n22104, QN => n26193);
   REGISTERS_reg_27_39_inst : DFF_X1 port map( D => n6128, CK => CLK, Q => 
                           n22103, QN => n26194);
   REGISTERS_reg_27_38_inst : DFF_X1 port map( D => n6127, CK => CLK, Q => 
                           n22102, QN => n26195);
   REGISTERS_reg_26_59_inst : DFF_X1 port map( D => n6212, CK => CLK, Q => 
                           n9312, QN => n26108);
   REGISTERS_reg_26_58_inst : DFF_X1 port map( D => n6211, CK => CLK, Q => 
                           n9317, QN => n26109);
   REGISTERS_reg_26_57_inst : DFF_X1 port map( D => n6210, CK => CLK, Q => 
                           n9322, QN => n26110);
   REGISTERS_reg_26_56_inst : DFF_X1 port map( D => n6209, CK => CLK, Q => 
                           n9327, QN => n26111);
   REGISTERS_reg_26_55_inst : DFF_X1 port map( D => n6208, CK => CLK, Q => 
                           n9332, QN => n26112);
   REGISTERS_reg_26_54_inst : DFF_X1 port map( D => n6207, CK => CLK, Q => 
                           n9337, QN => n26113);
   REGISTERS_reg_26_53_inst : DFF_X1 port map( D => n6206, CK => CLK, Q => 
                           n9342, QN => n26114);
   REGISTERS_reg_26_52_inst : DFF_X1 port map( D => n6205, CK => CLK, Q => 
                           n9347, QN => n26115);
   REGISTERS_reg_26_51_inst : DFF_X1 port map( D => n6204, CK => CLK, Q => 
                           n9352, QN => n26116);
   REGISTERS_reg_26_50_inst : DFF_X1 port map( D => n6203, CK => CLK, Q => 
                           n9357, QN => n26117);
   REGISTERS_reg_26_49_inst : DFF_X1 port map( D => n6202, CK => CLK, Q => 
                           n9362, QN => n26118);
   REGISTERS_reg_26_48_inst : DFF_X1 port map( D => n6201, CK => CLK, Q => 
                           n9367, QN => n26119);
   REGISTERS_reg_26_47_inst : DFF_X1 port map( D => n6200, CK => CLK, Q => 
                           n9372, QN => n26120);
   REGISTERS_reg_26_46_inst : DFF_X1 port map( D => n6199, CK => CLK, Q => 
                           n9377, QN => n26121);
   REGISTERS_reg_26_45_inst : DFF_X1 port map( D => n6198, CK => CLK, Q => 
                           n9382, QN => n26122);
   REGISTERS_reg_26_44_inst : DFF_X1 port map( D => n6197, CK => CLK, Q => 
                           n9387, QN => n26123);
   REGISTERS_reg_26_43_inst : DFF_X1 port map( D => n6196, CK => CLK, Q => 
                           n9392, QN => n26124);
   REGISTERS_reg_26_42_inst : DFF_X1 port map( D => n6195, CK => CLK, Q => 
                           n9397, QN => n26125);
   REGISTERS_reg_26_41_inst : DFF_X1 port map( D => n6194, CK => CLK, Q => 
                           n9402, QN => n26126);
   REGISTERS_reg_26_40_inst : DFF_X1 port map( D => n6193, CK => CLK, Q => 
                           n9407, QN => n26127);
   REGISTERS_reg_26_39_inst : DFF_X1 port map( D => n6192, CK => CLK, Q => 
                           n9412, QN => n26128);
   REGISTERS_reg_26_38_inst : DFF_X1 port map( D => n6191, CK => CLK, Q => 
                           n9417, QN => n26129);
   REGISTERS_reg_27_37_inst : DFF_X1 port map( D => n6126, CK => CLK, Q => 
                           n22101, QN => n26196);
   REGISTERS_reg_27_36_inst : DFF_X1 port map( D => n6125, CK => CLK, Q => 
                           n22100, QN => n26197);
   REGISTERS_reg_27_35_inst : DFF_X1 port map( D => n6124, CK => CLK, Q => 
                           n22099, QN => n26198);
   REGISTERS_reg_27_34_inst : DFF_X1 port map( D => n6123, CK => CLK, Q => 
                           n22098, QN => n26199);
   REGISTERS_reg_27_33_inst : DFF_X1 port map( D => n6122, CK => CLK, Q => 
                           n22097, QN => n26200);
   REGISTERS_reg_27_32_inst : DFF_X1 port map( D => n6121, CK => CLK, Q => 
                           n22096, QN => n26201);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n6120, CK => CLK, Q => 
                           n22095, QN => n26202);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n6119, CK => CLK, Q => 
                           n22094, QN => n26203);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n6118, CK => CLK, Q => 
                           n22093, QN => n26204);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n6117, CK => CLK, Q => 
                           n22092, QN => n26205);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n6116, CK => CLK, Q => 
                           n22091, QN => n26206);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n6115, CK => CLK, Q => 
                           n22090, QN => n26207);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n6114, CK => CLK, Q => 
                           n22089, QN => n26208);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n6113, CK => CLK, Q => 
                           n22088, QN => n26209);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n6112, CK => CLK, Q => 
                           n22087, QN => n26210);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n6111, CK => CLK, Q => 
                           n22086, QN => n26211);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n6110, CK => CLK, Q => 
                           n22085, QN => n26212);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n6109, CK => CLK, Q => 
                           n22084, QN => n26213);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n6108, CK => CLK, Q => 
                           n22083, QN => n26214);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n6107, CK => CLK, Q => 
                           n22082, QN => n26215);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n6106, CK => CLK, Q => 
                           n22081, QN => n26216);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n6105, CK => CLK, Q => 
                           n22080, QN => n26217);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n6104, CK => CLK, Q => 
                           n22079, QN => n26218);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n6103, CK => CLK, Q => 
                           n22078, QN => n26219);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n6102, CK => CLK, Q => 
                           n22077, QN => n26220);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n6101, CK => CLK, Q => 
                           n22076, QN => n26221);
   REGISTERS_reg_26_37_inst : DFF_X1 port map( D => n6190, CK => CLK, Q => 
                           n9422, QN => n26130);
   REGISTERS_reg_26_36_inst : DFF_X1 port map( D => n6189, CK => CLK, Q => 
                           n9427, QN => n26131);
   REGISTERS_reg_26_35_inst : DFF_X1 port map( D => n6188, CK => CLK, Q => 
                           n9432, QN => n26132);
   REGISTERS_reg_26_34_inst : DFF_X1 port map( D => n6187, CK => CLK, Q => 
                           n9437, QN => n26133);
   REGISTERS_reg_26_33_inst : DFF_X1 port map( D => n6186, CK => CLK, Q => 
                           n9442, QN => n26134);
   REGISTERS_reg_26_32_inst : DFF_X1 port map( D => n6185, CK => CLK, Q => 
                           n9447, QN => n26135);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n6184, CK => CLK, Q => 
                           n9452, QN => n26136);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n6183, CK => CLK, Q => 
                           n9457, QN => n26137);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n6182, CK => CLK, Q => 
                           n9462, QN => n26138);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n6181, CK => CLK, Q => 
                           n9467, QN => n26139);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n6180, CK => CLK, Q => 
                           n9472, QN => n26140);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n6179, CK => CLK, Q => 
                           n9477, QN => n26141);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n6178, CK => CLK, Q => 
                           n9482, QN => n26142);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n6177, CK => CLK, Q => 
                           n9487, QN => n26143);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n6176, CK => CLK, Q => 
                           n9492, QN => n26144);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n6175, CK => CLK, Q => 
                           n9497, QN => n26145);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n6174, CK => CLK, Q => 
                           n9502, QN => n26146);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n6173, CK => CLK, Q => 
                           n9507, QN => n26147);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n6172, CK => CLK, Q => 
                           n9512, QN => n26148);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n6171, CK => CLK, Q => 
                           n9517, QN => n26149);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n6170, CK => CLK, Q => 
                           n9522, QN => n26150);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n6169, CK => CLK, Q => 
                           n9527, QN => n26151);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n6168, CK => CLK, Q => 
                           n9532, QN => n26152);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n6167, CK => CLK, Q => 
                           n9537, QN => n26153);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n6166, CK => CLK, Q => 
                           n9542, QN => n26154);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n6165, CK => CLK, Q => 
                           n9547, QN => n26155);
   REGISTERS_reg_21_59_inst : DFF_X1 port map( D => n6532, CK => CLK, Q => 
                           n29956, QN => n26029);
   REGISTERS_reg_21_58_inst : DFF_X1 port map( D => n6531, CK => CLK, Q => 
                           n29955, QN => n26030);
   REGISTERS_reg_21_57_inst : DFF_X1 port map( D => n6530, CK => CLK, Q => 
                           n29954, QN => n26031);
   REGISTERS_reg_21_56_inst : DFF_X1 port map( D => n6529, CK => CLK, Q => 
                           n29953, QN => n26032);
   REGISTERS_reg_21_55_inst : DFF_X1 port map( D => n6528, CK => CLK, Q => 
                           n29952, QN => n26033);
   REGISTERS_reg_21_54_inst : DFF_X1 port map( D => n6527, CK => CLK, Q => 
                           n29951, QN => n26034);
   REGISTERS_reg_21_53_inst : DFF_X1 port map( D => n6526, CK => CLK, Q => 
                           n29950, QN => n26035);
   REGISTERS_reg_21_52_inst : DFF_X1 port map( D => n6525, CK => CLK, Q => 
                           n29949, QN => n26036);
   REGISTERS_reg_21_51_inst : DFF_X1 port map( D => n6524, CK => CLK, Q => 
                           n29948, QN => n26037);
   REGISTERS_reg_21_50_inst : DFF_X1 port map( D => n6523, CK => CLK, Q => 
                           n29947, QN => n26038);
   REGISTERS_reg_21_49_inst : DFF_X1 port map( D => n6522, CK => CLK, Q => 
                           n29946, QN => n26039);
   REGISTERS_reg_21_48_inst : DFF_X1 port map( D => n6521, CK => CLK, Q => 
                           n29945, QN => n26040);
   REGISTERS_reg_21_47_inst : DFF_X1 port map( D => n6520, CK => CLK, Q => 
                           n29944, QN => n26041);
   REGISTERS_reg_21_46_inst : DFF_X1 port map( D => n6519, CK => CLK, Q => 
                           n29943, QN => n26042);
   REGISTERS_reg_21_45_inst : DFF_X1 port map( D => n6518, CK => CLK, Q => 
                           n29942, QN => n26043);
   REGISTERS_reg_21_44_inst : DFF_X1 port map( D => n6517, CK => CLK, Q => 
                           n29941, QN => n26044);
   REGISTERS_reg_21_43_inst : DFF_X1 port map( D => n6516, CK => CLK, Q => 
                           n29940, QN => n26045);
   REGISTERS_reg_21_42_inst : DFF_X1 port map( D => n6515, CK => CLK, Q => 
                           n29939, QN => n26046);
   REGISTERS_reg_21_41_inst : DFF_X1 port map( D => n6514, CK => CLK, Q => 
                           n29938, QN => n26047);
   REGISTERS_reg_21_40_inst : DFF_X1 port map( D => n6513, CK => CLK, Q => 
                           n29937, QN => n26048);
   REGISTERS_reg_21_39_inst : DFF_X1 port map( D => n6512, CK => CLK, Q => 
                           n29936, QN => n26049);
   REGISTERS_reg_21_38_inst : DFF_X1 port map( D => n6511, CK => CLK, Q => 
                           n29935, QN => n26050);
   REGISTERS_reg_21_37_inst : DFF_X1 port map( D => n6510, CK => CLK, Q => 
                           n29934, QN => n26051);
   REGISTERS_reg_21_36_inst : DFF_X1 port map( D => n6509, CK => CLK, Q => 
                           n29933, QN => n26052);
   REGISTERS_reg_21_35_inst : DFF_X1 port map( D => n6508, CK => CLK, Q => 
                           n29932, QN => n26053);
   REGISTERS_reg_21_34_inst : DFF_X1 port map( D => n6507, CK => CLK, Q => 
                           n29931, QN => n26054);
   REGISTERS_reg_21_33_inst : DFF_X1 port map( D => n6506, CK => CLK, Q => 
                           n29930, QN => n26055);
   REGISTERS_reg_21_32_inst : DFF_X1 port map( D => n6505, CK => CLK, Q => 
                           n29929, QN => n26056);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n6504, CK => CLK, Q => 
                           n29928, QN => n26057);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n6503, CK => CLK, Q => 
                           n29927, QN => n26058);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n6502, CK => CLK, Q => 
                           n29926, QN => n26059);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n6501, CK => CLK, Q => 
                           n29925, QN => n26060);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n6500, CK => CLK, Q => 
                           n29924, QN => n26061);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n6499, CK => CLK, Q => 
                           n29923, QN => n26062);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n6498, CK => CLK, Q => 
                           n29922, QN => n26063);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n6497, CK => CLK, Q => 
                           n29921, QN => n26064);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n6496, CK => CLK, Q => 
                           n29920, QN => n26065);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n6495, CK => CLK, Q => 
                           n29919, QN => n26066);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n6494, CK => CLK, Q => 
                           n29918, QN => n26067);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n6493, CK => CLK, Q => 
                           n29917, QN => n26068);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n6492, CK => CLK, Q => 
                           n29916, QN => n26069);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n6491, CK => CLK, Q => 
                           n29915, QN => n26070);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n6490, CK => CLK, Q => 
                           n29914, QN => n26071);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n6489, CK => CLK, Q => 
                           n29913, QN => n26072);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n6488, CK => CLK, Q => 
                           n29912, QN => n26073);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n6487, CK => CLK, Q => 
                           n29911, QN => n26074);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n6486, CK => CLK, Q => 
                           n29910, QN => n26075);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n6485, CK => CLK, Q => 
                           n29909, QN => n26076);
   REGISTERS_reg_20_59_inst : DFF_X1 port map( D => n6596, CK => CLK, Q => 
                           n29908, QN => n25963);
   REGISTERS_reg_20_58_inst : DFF_X1 port map( D => n6595, CK => CLK, Q => 
                           n29907, QN => n25964);
   REGISTERS_reg_20_57_inst : DFF_X1 port map( D => n6594, CK => CLK, Q => 
                           n29906, QN => n25965);
   REGISTERS_reg_20_56_inst : DFF_X1 port map( D => n6593, CK => CLK, Q => 
                           n29905, QN => n25966);
   REGISTERS_reg_20_55_inst : DFF_X1 port map( D => n6592, CK => CLK, Q => 
                           n29904, QN => n25967);
   REGISTERS_reg_20_54_inst : DFF_X1 port map( D => n6591, CK => CLK, Q => 
                           n29903, QN => n25968);
   REGISTERS_reg_20_53_inst : DFF_X1 port map( D => n6590, CK => CLK, Q => 
                           n29902, QN => n25969);
   REGISTERS_reg_20_52_inst : DFF_X1 port map( D => n6589, CK => CLK, Q => 
                           n29901, QN => n25970);
   REGISTERS_reg_20_51_inst : DFF_X1 port map( D => n6588, CK => CLK, Q => 
                           n29900, QN => n25971);
   REGISTERS_reg_20_50_inst : DFF_X1 port map( D => n6587, CK => CLK, Q => 
                           n29899, QN => n25972);
   REGISTERS_reg_20_49_inst : DFF_X1 port map( D => n6586, CK => CLK, Q => 
                           n29898, QN => n25973);
   REGISTERS_reg_20_48_inst : DFF_X1 port map( D => n6585, CK => CLK, Q => 
                           n29897, QN => n25974);
   REGISTERS_reg_20_47_inst : DFF_X1 port map( D => n6584, CK => CLK, Q => 
                           n29896, QN => n25975);
   REGISTERS_reg_20_46_inst : DFF_X1 port map( D => n6583, CK => CLK, Q => 
                           n29895, QN => n25976);
   REGISTERS_reg_20_45_inst : DFF_X1 port map( D => n6582, CK => CLK, Q => 
                           n29894, QN => n25977);
   REGISTERS_reg_20_44_inst : DFF_X1 port map( D => n6581, CK => CLK, Q => 
                           n29893, QN => n25978);
   REGISTERS_reg_20_43_inst : DFF_X1 port map( D => n6580, CK => CLK, Q => 
                           n29892, QN => n25979);
   REGISTERS_reg_20_42_inst : DFF_X1 port map( D => n6579, CK => CLK, Q => 
                           n29891, QN => n25980);
   REGISTERS_reg_20_41_inst : DFF_X1 port map( D => n6578, CK => CLK, Q => 
                           n29890, QN => n25981);
   REGISTERS_reg_20_40_inst : DFF_X1 port map( D => n6577, CK => CLK, Q => 
                           n29889, QN => n25982);
   REGISTERS_reg_20_39_inst : DFF_X1 port map( D => n6576, CK => CLK, Q => 
                           n29888, QN => n25983);
   REGISTERS_reg_20_38_inst : DFF_X1 port map( D => n6575, CK => CLK, Q => 
                           n29887, QN => n25984);
   REGISTERS_reg_20_37_inst : DFF_X1 port map( D => n6574, CK => CLK, Q => 
                           n29886, QN => n25985);
   REGISTERS_reg_20_36_inst : DFF_X1 port map( D => n6573, CK => CLK, Q => 
                           n29885, QN => n25986);
   REGISTERS_reg_20_35_inst : DFF_X1 port map( D => n6572, CK => CLK, Q => 
                           n29884, QN => n25987);
   REGISTERS_reg_20_34_inst : DFF_X1 port map( D => n6571, CK => CLK, Q => 
                           n29883, QN => n25988);
   REGISTERS_reg_20_33_inst : DFF_X1 port map( D => n6570, CK => CLK, Q => 
                           n29882, QN => n25989);
   REGISTERS_reg_20_32_inst : DFF_X1 port map( D => n6569, CK => CLK, Q => 
                           n29881, QN => n25990);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n6568, CK => CLK, Q => 
                           n29880, QN => n25991);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n6567, CK => CLK, Q => 
                           n29879, QN => n25992);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n6566, CK => CLK, Q => 
                           n29878, QN => n25993);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n6565, CK => CLK, Q => 
                           n29877, QN => n25994);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n6564, CK => CLK, Q => 
                           n29876, QN => n25995);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n6563, CK => CLK, Q => 
                           n29875, QN => n25996);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n6562, CK => CLK, Q => 
                           n29874, QN => n25997);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n6561, CK => CLK, Q => 
                           n29873, QN => n25998);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n6560, CK => CLK, Q => 
                           n29872, QN => n25999);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n6559, CK => CLK, Q => 
                           n29871, QN => n26000);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n6558, CK => CLK, Q => 
                           n29870, QN => n26001);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n6557, CK => CLK, Q => 
                           n29869, QN => n26002);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n6556, CK => CLK, Q => 
                           n29868, QN => n26003);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n6555, CK => CLK, Q => 
                           n29867, QN => n26004);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n6554, CK => CLK, Q => 
                           n29866, QN => n26005);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n6553, CK => CLK, Q => 
                           n29865, QN => n26006);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n6552, CK => CLK, Q => 
                           n29864, QN => n26007);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n6551, CK => CLK, Q => 
                           n29863, QN => n26008);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n6550, CK => CLK, Q => 
                           n29862, QN => n26009);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n6549, CK => CLK, Q => 
                           n29861, QN => n26010);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n6740, CK => CLK, Q => 
                           n21870, QN => n25928);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n6739, CK => CLK, Q => 
                           n21869, QN => n25929);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n6738, CK => CLK, Q => 
                           n21868, QN => n25930);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n6737, CK => CLK, Q => 
                           n21867, QN => n25931);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n6736, CK => CLK, Q => 
                           n21866, QN => n25932);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n6735, CK => CLK, Q => 
                           n21865, QN => n25933);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n6734, CK => CLK, Q => 
                           n21864, QN => n25934);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n6733, CK => CLK, Q => 
                           n21863, QN => n25935);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n6732, CK => CLK, Q => 
                           n21862, QN => n25936);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n6731, CK => CLK, Q => 
                           n21861, QN => n25937);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n6730, CK => CLK, Q => 
                           n21860, QN => n25938);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n6729, CK => CLK, Q => 
                           n21859, QN => n25939);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n6804, CK => CLK, Q => 
                           n9553, QN => n25861);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n6803, CK => CLK, Q => 
                           n9558, QN => n25862);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n6802, CK => CLK, Q => n9563
                           , QN => n25863);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n6801, CK => CLK, Q => n9568
                           , QN => n25864);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n6800, CK => CLK, Q => n9573
                           , QN => n25865);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n6799, CK => CLK, Q => n9578
                           , QN => n25866);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n6798, CK => CLK, Q => n9583
                           , QN => n25867);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n6797, CK => CLK, Q => n9588
                           , QN => n25868);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n6796, CK => CLK, Q => n9593
                           , QN => n25869);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n6795, CK => CLK, Q => n9598
                           , QN => n25870);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n6794, CK => CLK, Q => n9603
                           , QN => n25871);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n6793, CK => CLK, Q => n9608
                           , QN => n25872);
   REGISTERS_reg_17_59_inst : DFF_X1 port map( D => n6788, CK => CLK, Q => 
                           n21918, QN => n25880);
   REGISTERS_reg_17_58_inst : DFF_X1 port map( D => n6787, CK => CLK, Q => 
                           n21917, QN => n25881);
   REGISTERS_reg_17_57_inst : DFF_X1 port map( D => n6786, CK => CLK, Q => 
                           n21916, QN => n25882);
   REGISTERS_reg_17_56_inst : DFF_X1 port map( D => n6785, CK => CLK, Q => 
                           n21915, QN => n25883);
   REGISTERS_reg_17_55_inst : DFF_X1 port map( D => n6784, CK => CLK, Q => 
                           n21914, QN => n25884);
   REGISTERS_reg_17_54_inst : DFF_X1 port map( D => n6783, CK => CLK, Q => 
                           n21913, QN => n25885);
   REGISTERS_reg_17_53_inst : DFF_X1 port map( D => n6782, CK => CLK, Q => 
                           n21912, QN => n25886);
   REGISTERS_reg_17_52_inst : DFF_X1 port map( D => n6781, CK => CLK, Q => 
                           n21911, QN => n25887);
   REGISTERS_reg_17_51_inst : DFF_X1 port map( D => n6780, CK => CLK, Q => 
                           n21910, QN => n25888);
   REGISTERS_reg_17_50_inst : DFF_X1 port map( D => n6779, CK => CLK, Q => 
                           n21909, QN => n25889);
   REGISTERS_reg_17_49_inst : DFF_X1 port map( D => n6778, CK => CLK, Q => 
                           n21908, QN => n25890);
   REGISTERS_reg_17_48_inst : DFF_X1 port map( D => n6777, CK => CLK, Q => 
                           n21907, QN => n25891);
   REGISTERS_reg_17_47_inst : DFF_X1 port map( D => n6776, CK => CLK, Q => 
                           n21906, QN => n25892);
   REGISTERS_reg_17_46_inst : DFF_X1 port map( D => n6775, CK => CLK, Q => 
                           n21905, QN => n25893);
   REGISTERS_reg_17_45_inst : DFF_X1 port map( D => n6774, CK => CLK, Q => 
                           n21904, QN => n25894);
   REGISTERS_reg_17_44_inst : DFF_X1 port map( D => n6773, CK => CLK, Q => 
                           n21903, QN => n25895);
   REGISTERS_reg_17_43_inst : DFF_X1 port map( D => n6772, CK => CLK, Q => 
                           n21902, QN => n25896);
   REGISTERS_reg_17_42_inst : DFF_X1 port map( D => n6771, CK => CLK, Q => 
                           n21901, QN => n25897);
   REGISTERS_reg_17_41_inst : DFF_X1 port map( D => n6770, CK => CLK, Q => 
                           n21900, QN => n25898);
   REGISTERS_reg_17_40_inst : DFF_X1 port map( D => n6769, CK => CLK, Q => 
                           n21899, QN => n25899);
   REGISTERS_reg_17_39_inst : DFF_X1 port map( D => n6768, CK => CLK, Q => 
                           n21898, QN => n25900);
   REGISTERS_reg_17_38_inst : DFF_X1 port map( D => n6767, CK => CLK, Q => 
                           n21897, QN => n25901);
   REGISTERS_reg_16_59_inst : DFF_X1 port map( D => n6852, CK => CLK, Q => 
                           n9313, QN => n25813);
   REGISTERS_reg_16_58_inst : DFF_X1 port map( D => n6851, CK => CLK, Q => 
                           n9318, QN => n25814);
   REGISTERS_reg_16_57_inst : DFF_X1 port map( D => n6850, CK => CLK, Q => 
                           n9323, QN => n25815);
   REGISTERS_reg_16_56_inst : DFF_X1 port map( D => n6849, CK => CLK, Q => 
                           n9328, QN => n25816);
   REGISTERS_reg_16_55_inst : DFF_X1 port map( D => n6848, CK => CLK, Q => 
                           n9333, QN => n25817);
   REGISTERS_reg_16_54_inst : DFF_X1 port map( D => n6847, CK => CLK, Q => 
                           n9338, QN => n25818);
   REGISTERS_reg_16_53_inst : DFF_X1 port map( D => n6846, CK => CLK, Q => 
                           n9343, QN => n25819);
   REGISTERS_reg_16_52_inst : DFF_X1 port map( D => n6845, CK => CLK, Q => 
                           n9348, QN => n25820);
   REGISTERS_reg_16_51_inst : DFF_X1 port map( D => n6844, CK => CLK, Q => 
                           n9353, QN => n25821);
   REGISTERS_reg_16_50_inst : DFF_X1 port map( D => n6843, CK => CLK, Q => 
                           n9358, QN => n25822);
   REGISTERS_reg_16_49_inst : DFF_X1 port map( D => n6842, CK => CLK, Q => 
                           n9363, QN => n25823);
   REGISTERS_reg_16_48_inst : DFF_X1 port map( D => n6841, CK => CLK, Q => 
                           n9368, QN => n25824);
   REGISTERS_reg_16_47_inst : DFF_X1 port map( D => n6840, CK => CLK, Q => 
                           n9373, QN => n25825);
   REGISTERS_reg_16_46_inst : DFF_X1 port map( D => n6839, CK => CLK, Q => 
                           n9378, QN => n25826);
   REGISTERS_reg_16_45_inst : DFF_X1 port map( D => n6838, CK => CLK, Q => 
                           n9383, QN => n25827);
   REGISTERS_reg_16_44_inst : DFF_X1 port map( D => n6837, CK => CLK, Q => 
                           n9388, QN => n25828);
   REGISTERS_reg_16_43_inst : DFF_X1 port map( D => n6836, CK => CLK, Q => 
                           n9393, QN => n25829);
   REGISTERS_reg_16_42_inst : DFF_X1 port map( D => n6835, CK => CLK, Q => 
                           n9398, QN => n25830);
   REGISTERS_reg_16_41_inst : DFF_X1 port map( D => n6834, CK => CLK, Q => 
                           n9403, QN => n25831);
   REGISTERS_reg_16_40_inst : DFF_X1 port map( D => n6833, CK => CLK, Q => 
                           n9408, QN => n25832);
   REGISTERS_reg_16_39_inst : DFF_X1 port map( D => n6832, CK => CLK, Q => 
                           n9413, QN => n25833);
   REGISTERS_reg_16_38_inst : DFF_X1 port map( D => n6831, CK => CLK, Q => 
                           n9418, QN => n25834);
   REGISTERS_reg_17_37_inst : DFF_X1 port map( D => n6766, CK => CLK, Q => 
                           n21896, QN => n25902);
   REGISTERS_reg_17_36_inst : DFF_X1 port map( D => n6765, CK => CLK, Q => 
                           n21895, QN => n25903);
   REGISTERS_reg_17_35_inst : DFF_X1 port map( D => n6764, CK => CLK, Q => 
                           n21894, QN => n25904);
   REGISTERS_reg_17_34_inst : DFF_X1 port map( D => n6763, CK => CLK, Q => 
                           n21893, QN => n25905);
   REGISTERS_reg_17_33_inst : DFF_X1 port map( D => n6762, CK => CLK, Q => 
                           n21892, QN => n25906);
   REGISTERS_reg_17_32_inst : DFF_X1 port map( D => n6761, CK => CLK, Q => 
                           n21891, QN => n25907);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n6760, CK => CLK, Q => 
                           n21890, QN => n25908);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n6759, CK => CLK, Q => 
                           n21889, QN => n25909);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n6758, CK => CLK, Q => 
                           n21888, QN => n25910);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n6757, CK => CLK, Q => 
                           n21887, QN => n25911);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n6756, CK => CLK, Q => 
                           n21886, QN => n25912);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n6755, CK => CLK, Q => 
                           n21885, QN => n25913);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n6754, CK => CLK, Q => 
                           n21884, QN => n25914);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n6753, CK => CLK, Q => 
                           n21883, QN => n25915);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n6752, CK => CLK, Q => 
                           n21882, QN => n25916);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n6751, CK => CLK, Q => 
                           n21881, QN => n25917);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n6750, CK => CLK, Q => 
                           n21880, QN => n25918);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n6749, CK => CLK, Q => 
                           n21879, QN => n25919);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n6748, CK => CLK, Q => 
                           n21878, QN => n25920);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n6747, CK => CLK, Q => 
                           n21877, QN => n25921);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n6746, CK => CLK, Q => 
                           n21876, QN => n25922);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n6745, CK => CLK, Q => 
                           n21875, QN => n25923);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n6744, CK => CLK, Q => 
                           n21874, QN => n25924);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n6743, CK => CLK, Q => 
                           n21873, QN => n25925);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n6742, CK => CLK, Q => 
                           n21872, QN => n25926);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n6741, CK => CLK, Q => 
                           n21871, QN => n25927);
   REGISTERS_reg_16_37_inst : DFF_X1 port map( D => n6830, CK => CLK, Q => 
                           n9423, QN => n25835);
   REGISTERS_reg_16_36_inst : DFF_X1 port map( D => n6829, CK => CLK, Q => 
                           n9428, QN => n25836);
   REGISTERS_reg_16_35_inst : DFF_X1 port map( D => n6828, CK => CLK, Q => 
                           n9433, QN => n25837);
   REGISTERS_reg_16_34_inst : DFF_X1 port map( D => n6827, CK => CLK, Q => 
                           n9438, QN => n25838);
   REGISTERS_reg_16_33_inst : DFF_X1 port map( D => n6826, CK => CLK, Q => 
                           n9443, QN => n25839);
   REGISTERS_reg_16_32_inst : DFF_X1 port map( D => n6825, CK => CLK, Q => 
                           n9448, QN => n25840);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n6824, CK => CLK, Q => 
                           n9453, QN => n25841);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n6823, CK => CLK, Q => 
                           n9458, QN => n25842);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n6822, CK => CLK, Q => 
                           n9463, QN => n25843);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n6821, CK => CLK, Q => 
                           n9468, QN => n25844);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n6820, CK => CLK, Q => 
                           n9473, QN => n25845);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n6819, CK => CLK, Q => 
                           n9478, QN => n25846);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n6818, CK => CLK, Q => 
                           n9483, QN => n25847);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n6817, CK => CLK, Q => 
                           n9488, QN => n25848);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n6816, CK => CLK, Q => 
                           n9493, QN => n25849);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n6815, CK => CLK, Q => 
                           n9498, QN => n25850);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n6814, CK => CLK, Q => 
                           n9503, QN => n25851);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n6813, CK => CLK, Q => 
                           n9508, QN => n25852);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n6812, CK => CLK, Q => 
                           n9513, QN => n25853);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n6811, CK => CLK, Q => 
                           n9518, QN => n25854);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n6810, CK => CLK, Q => 
                           n9523, QN => n25855);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n6809, CK => CLK, Q => 
                           n9528, QN => n25856);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n6808, CK => CLK, Q => 
                           n9533, QN => n25857);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n6807, CK => CLK, Q => 
                           n9538, QN => n25858);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n6806, CK => CLK, Q => 
                           n9543, QN => n25859);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n6805, CK => CLK, Q => 
                           n9548, QN => n25860);
   REGISTERS_reg_6_63_inst : DFF_X1 port map( D => n7496, CK => CLK, Q => n9290
                           , QN => n25386);
   REGISTERS_reg_6_62_inst : DFF_X1 port map( D => n7495, CK => CLK, Q => n9295
                           , QN => n25388);
   REGISTERS_reg_6_61_inst : DFF_X1 port map( D => n7494, CK => CLK, Q => n9300
                           , QN => n25389);
   REGISTERS_reg_6_60_inst : DFF_X1 port map( D => n7493, CK => CLK, Q => n9305
                           , QN => n25390);
   REGISTERS_reg_2_63_inst : DFF_X1 port map( D => n7752, CK => CLK, Q => n9289
                           , QN => n25237);
   REGISTERS_reg_2_62_inst : DFF_X1 port map( D => n7751, CK => CLK, Q => n9294
                           , QN => n25239);
   REGISTERS_reg_2_61_inst : DFF_X1 port map( D => n7750, CK => CLK, Q => n9299
                           , QN => n25240);
   REGISTERS_reg_2_60_inst : DFF_X1 port map( D => n7749, CK => CLK, Q => n9304
                           , QN => n25241);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n7827, CK => CLK, Q => 
                           n29860, QN => n25209);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n7826, CK => CLK, Q => n29859
                           , QN => n25211);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n7825, CK => CLK, Q => n29858
                           , QN => n25213);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n7824, CK => CLK, Q => n29857
                           , QN => n25215);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n7823, CK => CLK, Q => n29856
                           , QN => n25217);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n7822, CK => CLK, Q => n29855
                           , QN => n25219);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n7821, CK => CLK, Q => n29854
                           , QN => n25221);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n7820, CK => CLK, Q => n29853
                           , QN => n25223);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n7819, CK => CLK, Q => n29852
                           , QN => n25225);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n7818, CK => CLK, Q => n29851
                           , QN => n25227);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n7817, CK => CLK, Q => n29850
                           , QN => n25229);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n7571, CK => CLK, Q => 
                           n29849, QN => n25371);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n7570, CK => CLK, Q => n29848
                           , QN => n25372);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n7569, CK => CLK, Q => n29847
                           , QN => n25373);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n7568, CK => CLK, Q => n29846
                           , QN => n25374);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n7567, CK => CLK, Q => n29845
                           , QN => n25375);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n7566, CK => CLK, Q => n29844
                           , QN => n25376);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n7565, CK => CLK, Q => n29843
                           , QN => n25377);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n7564, CK => CLK, Q => n29842
                           , QN => n25378);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n7563, CK => CLK, Q => n29841
                           , QN => n25379);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n7562, CK => CLK, Q => n29840
                           , QN => n25380);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n7561, CK => CLK, Q => n29839
                           , QN => n25381);
   REGISTERS_reg_13_63_inst : DFF_X1 port map( D => n7048, CK => CLK, Q => 
                           n22242, QN => n25737);
   REGISTERS_reg_13_62_inst : DFF_X1 port map( D => n7047, CK => CLK, Q => 
                           n22241, QN => n25739);
   REGISTERS_reg_13_61_inst : DFF_X1 port map( D => n7046, CK => CLK, Q => 
                           n22240, QN => n25740);
   REGISTERS_reg_13_60_inst : DFF_X1 port map( D => n7045, CK => CLK, Q => 
                           n22239, QN => n25741);
   REGISTERS_reg_9_63_inst : DFF_X1 port map( D => n7304, CK => CLK, Q => 
                           n22015, QN => n25589);
   REGISTERS_reg_9_62_inst : DFF_X1 port map( D => n7303, CK => CLK, Q => 
                           n22014, QN => n25591);
   REGISTERS_reg_9_61_inst : DFF_X1 port map( D => n7302, CK => CLK, Q => 
                           n22013, QN => n25592);
   REGISTERS_reg_9_60_inst : DFF_X1 port map( D => n7301, CK => CLK, Q => 
                           n22012, QN => n25593);
   REGISTERS_reg_7_63_inst : DFF_X1 port map( D => n7432, CK => CLK, Q => 
                           n21926, QN => n25456);
   REGISTERS_reg_7_62_inst : DFF_X1 port map( D => n7431, CK => CLK, Q => 
                           n21925, QN => n25458);
   REGISTERS_reg_7_61_inst : DFF_X1 port map( D => n7430, CK => CLK, Q => 
                           n21924, QN => n25459);
   REGISTERS_reg_7_60_inst : DFF_X1 port map( D => n7429, CK => CLK, Q => 
                           n21923, QN => n25460);
   REGISTERS_reg_3_63_inst : DFF_X1 port map( D => n7688, CK => CLK, Q => 
                           n21858, QN => n25304);
   REGISTERS_reg_3_62_inst : DFF_X1 port map( D => n7687, CK => CLK, Q => 
                           n21857, QN => n25306);
   REGISTERS_reg_3_61_inst : DFF_X1 port map( D => n7686, CK => CLK, Q => 
                           n21856, QN => n25307);
   REGISTERS_reg_3_60_inst : DFF_X1 port map( D => n7685, CK => CLK, Q => 
                           n21855, QN => n25308);
   REGISTERS_reg_12_63_inst : DFF_X1 port map( D => n7112, CK => CLK, Q => 
                           n9673, QN => n25671);
   REGISTERS_reg_12_62_inst : DFF_X1 port map( D => n7111, CK => CLK, Q => 
                           n9674, QN => n25673);
   REGISTERS_reg_12_61_inst : DFF_X1 port map( D => n7110, CK => CLK, Q => 
                           n9675, QN => n25674);
   REGISTERS_reg_12_60_inst : DFF_X1 port map( D => n7109, CK => CLK, Q => 
                           n9676, QN => n25675);
   REGISTERS_reg_8_63_inst : DFF_X1 port map( D => n7368, CK => CLK, Q => n9291
                           , QN => n25522);
   REGISTERS_reg_8_62_inst : DFF_X1 port map( D => n7367, CK => CLK, Q => n9296
                           , QN => n25524);
   REGISTERS_reg_8_61_inst : DFF_X1 port map( D => n7366, CK => CLK, Q => n9301
                           , QN => n25525);
   REGISTERS_reg_8_60_inst : DFF_X1 port map( D => n7365, CK => CLK, Q => n9306
                           , QN => n25526);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n7187, CK => CLK, Q => 
                           n29838, QN => n25657);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n7186, CK => CLK, Q => 
                           n29837, QN => n25658);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n7185, CK => CLK, Q => 
                           n29836, QN => n25659);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n7184, CK => CLK, Q => 
                           n29835, QN => n25660);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n7183, CK => CLK, Q => 
                           n29834, QN => n25661);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n7182, CK => CLK, Q => 
                           n29833, QN => n25662);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n7181, CK => CLK, Q => 
                           n29832, QN => n25663);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n7180, CK => CLK, Q => 
                           n29831, QN => n25664);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n7179, CK => CLK, Q => 
                           n29830, QN => n25665);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n7178, CK => CLK, Q => 
                           n29829, QN => n25666);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n7177, CK => CLK, Q => 
                           n29828, QN => n25667);
   REGISTERS_reg_6_59_inst : DFF_X1 port map( D => n7492, CK => CLK, Q => n9310
                           , QN => n25391);
   REGISTERS_reg_6_58_inst : DFF_X1 port map( D => n7491, CK => CLK, Q => n9315
                           , QN => n25392);
   REGISTERS_reg_6_57_inst : DFF_X1 port map( D => n7490, CK => CLK, Q => n9320
                           , QN => n25393);
   REGISTERS_reg_6_56_inst : DFF_X1 port map( D => n7489, CK => CLK, Q => n9325
                           , QN => n25394);
   REGISTERS_reg_6_55_inst : DFF_X1 port map( D => n7488, CK => CLK, Q => n9330
                           , QN => n25395);
   REGISTERS_reg_6_54_inst : DFF_X1 port map( D => n7487, CK => CLK, Q => n9335
                           , QN => n25396);
   REGISTERS_reg_6_53_inst : DFF_X1 port map( D => n7486, CK => CLK, Q => n9340
                           , QN => n25397);
   REGISTERS_reg_6_52_inst : DFF_X1 port map( D => n7485, CK => CLK, Q => n9345
                           , QN => n25398);
   REGISTERS_reg_6_51_inst : DFF_X1 port map( D => n7484, CK => CLK, Q => n9350
                           , QN => n25399);
   REGISTERS_reg_6_50_inst : DFF_X1 port map( D => n7483, CK => CLK, Q => n9355
                           , QN => n25400);
   REGISTERS_reg_6_49_inst : DFF_X1 port map( D => n7482, CK => CLK, Q => n9360
                           , QN => n25401);
   REGISTERS_reg_6_48_inst : DFF_X1 port map( D => n7481, CK => CLK, Q => n9365
                           , QN => n25402);
   REGISTERS_reg_6_47_inst : DFF_X1 port map( D => n7480, CK => CLK, Q => n9370
                           , QN => n25403);
   REGISTERS_reg_6_46_inst : DFF_X1 port map( D => n7479, CK => CLK, Q => n9375
                           , QN => n25404);
   REGISTERS_reg_6_45_inst : DFF_X1 port map( D => n7478, CK => CLK, Q => n9380
                           , QN => n25405);
   REGISTERS_reg_6_44_inst : DFF_X1 port map( D => n7477, CK => CLK, Q => n9385
                           , QN => n25406);
   REGISTERS_reg_6_43_inst : DFF_X1 port map( D => n7476, CK => CLK, Q => n9390
                           , QN => n25407);
   REGISTERS_reg_6_42_inst : DFF_X1 port map( D => n7475, CK => CLK, Q => n9395
                           , QN => n25408);
   REGISTERS_reg_6_41_inst : DFF_X1 port map( D => n7474, CK => CLK, Q => n9400
                           , QN => n25409);
   REGISTERS_reg_6_40_inst : DFF_X1 port map( D => n7473, CK => CLK, Q => n9405
                           , QN => n25410);
   REGISTERS_reg_6_39_inst : DFF_X1 port map( D => n7472, CK => CLK, Q => n9410
                           , QN => n25411);
   REGISTERS_reg_6_38_inst : DFF_X1 port map( D => n7471, CK => CLK, Q => n9415
                           , QN => n25412);
   REGISTERS_reg_6_37_inst : DFF_X1 port map( D => n7470, CK => CLK, Q => n9420
                           , QN => n25413);
   REGISTERS_reg_6_36_inst : DFF_X1 port map( D => n7469, CK => CLK, Q => n9425
                           , QN => n25414);
   REGISTERS_reg_6_35_inst : DFF_X1 port map( D => n7468, CK => CLK, Q => n9430
                           , QN => n25415);
   REGISTERS_reg_6_34_inst : DFF_X1 port map( D => n7467, CK => CLK, Q => n9435
                           , QN => n25416);
   REGISTERS_reg_6_33_inst : DFF_X1 port map( D => n7466, CK => CLK, Q => n9440
                           , QN => n25417);
   REGISTERS_reg_6_32_inst : DFF_X1 port map( D => n7465, CK => CLK, Q => n9445
                           , QN => n25418);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n7464, CK => CLK, Q => n9450
                           , QN => n25419);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n7463, CK => CLK, Q => n9455
                           , QN => n25420);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n7462, CK => CLK, Q => n9460
                           , QN => n25421);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n7461, CK => CLK, Q => n9465
                           , QN => n25422);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n7460, CK => CLK, Q => n9470
                           , QN => n25423);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n7459, CK => CLK, Q => n9475
                           , QN => n25424);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n7458, CK => CLK, Q => n9480
                           , QN => n25425);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n7457, CK => CLK, Q => n9485
                           , QN => n25426);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n7456, CK => CLK, Q => n9490
                           , QN => n25427);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n7455, CK => CLK, Q => n9495
                           , QN => n25428);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n7454, CK => CLK, Q => n9500
                           , QN => n25429);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n7453, CK => CLK, Q => n9505
                           , QN => n25430);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n7452, CK => CLK, Q => n9510
                           , QN => n25431);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n7451, CK => CLK, Q => n9515
                           , QN => n25432);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n7450, CK => CLK, Q => n9520
                           , QN => n25433);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n7449, CK => CLK, Q => n9525
                           , QN => n25434);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n7448, CK => CLK, Q => n9530
                           , QN => n25435);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n7447, CK => CLK, Q => n9535
                           , QN => n25436);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n7446, CK => CLK, Q => n9540
                           , QN => n25437);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n7445, CK => CLK, Q => n9545
                           , QN => n25438);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n7444, CK => CLK, Q => n9550
                           , QN => n25439);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n7443, CK => CLK, Q => n9555
                           , QN => n25440);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n7442, CK => CLK, Q => n9560,
                           QN => n25441);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n7441, CK => CLK, Q => n9565,
                           QN => n25442);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n7440, CK => CLK, Q => n9570,
                           QN => n25443);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n7439, CK => CLK, Q => n9575,
                           QN => n25444);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n7438, CK => CLK, Q => n9580,
                           QN => n25445);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n7437, CK => CLK, Q => n9585,
                           QN => n25446);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n7436, CK => CLK, Q => n9590,
                           QN => n25447);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n7435, CK => CLK, Q => n9595,
                           QN => n25448);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n7434, CK => CLK, Q => n9600,
                           QN => n25449);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n7433, CK => CLK, Q => n9605,
                           QN => n25450);
   REGISTERS_reg_2_59_inst : DFF_X1 port map( D => n7748, CK => CLK, Q => n9309
                           , QN => n25242);
   REGISTERS_reg_2_58_inst : DFF_X1 port map( D => n7747, CK => CLK, Q => n9314
                           , QN => n25243);
   REGISTERS_reg_2_57_inst : DFF_X1 port map( D => n7746, CK => CLK, Q => n9319
                           , QN => n25244);
   REGISTERS_reg_2_56_inst : DFF_X1 port map( D => n7745, CK => CLK, Q => n9324
                           , QN => n25245);
   REGISTERS_reg_2_55_inst : DFF_X1 port map( D => n7744, CK => CLK, Q => n9329
                           , QN => n25246);
   REGISTERS_reg_2_54_inst : DFF_X1 port map( D => n7743, CK => CLK, Q => n9334
                           , QN => n25247);
   REGISTERS_reg_2_53_inst : DFF_X1 port map( D => n7742, CK => CLK, Q => n9339
                           , QN => n25248);
   REGISTERS_reg_2_52_inst : DFF_X1 port map( D => n7741, CK => CLK, Q => n9344
                           , QN => n25249);
   REGISTERS_reg_2_51_inst : DFF_X1 port map( D => n7740, CK => CLK, Q => n9349
                           , QN => n25250);
   REGISTERS_reg_2_50_inst : DFF_X1 port map( D => n7739, CK => CLK, Q => n9354
                           , QN => n25251);
   REGISTERS_reg_2_49_inst : DFF_X1 port map( D => n7738, CK => CLK, Q => n9359
                           , QN => n25252);
   REGISTERS_reg_2_48_inst : DFF_X1 port map( D => n7737, CK => CLK, Q => n9364
                           , QN => n25253);
   REGISTERS_reg_2_47_inst : DFF_X1 port map( D => n7736, CK => CLK, Q => n9369
                           , QN => n25254);
   REGISTERS_reg_2_46_inst : DFF_X1 port map( D => n7735, CK => CLK, Q => n9374
                           , QN => n25255);
   REGISTERS_reg_2_45_inst : DFF_X1 port map( D => n7734, CK => CLK, Q => n9379
                           , QN => n25256);
   REGISTERS_reg_2_44_inst : DFF_X1 port map( D => n7733, CK => CLK, Q => n9384
                           , QN => n25257);
   REGISTERS_reg_2_43_inst : DFF_X1 port map( D => n7732, CK => CLK, Q => n9389
                           , QN => n25258);
   REGISTERS_reg_2_42_inst : DFF_X1 port map( D => n7731, CK => CLK, Q => n9394
                           , QN => n25259);
   REGISTERS_reg_2_41_inst : DFF_X1 port map( D => n7730, CK => CLK, Q => n9399
                           , QN => n25260);
   REGISTERS_reg_2_40_inst : DFF_X1 port map( D => n7729, CK => CLK, Q => n9404
                           , QN => n25261);
   REGISTERS_reg_2_39_inst : DFF_X1 port map( D => n7728, CK => CLK, Q => n9409
                           , QN => n25262);
   REGISTERS_reg_2_38_inst : DFF_X1 port map( D => n7727, CK => CLK, Q => n9414
                           , QN => n25263);
   REGISTERS_reg_2_37_inst : DFF_X1 port map( D => n7726, CK => CLK, Q => n9419
                           , QN => n25264);
   REGISTERS_reg_2_36_inst : DFF_X1 port map( D => n7725, CK => CLK, Q => n9424
                           , QN => n25265);
   REGISTERS_reg_2_35_inst : DFF_X1 port map( D => n7724, CK => CLK, Q => n9429
                           , QN => n25266);
   REGISTERS_reg_2_34_inst : DFF_X1 port map( D => n7723, CK => CLK, Q => n9434
                           , QN => n25267);
   REGISTERS_reg_2_33_inst : DFF_X1 port map( D => n7722, CK => CLK, Q => n9439
                           , QN => n25268);
   REGISTERS_reg_2_32_inst : DFF_X1 port map( D => n7721, CK => CLK, Q => n9444
                           , QN => n25269);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n7720, CK => CLK, Q => n9449
                           , QN => n25270);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n7719, CK => CLK, Q => n9454
                           , QN => n25271);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n7718, CK => CLK, Q => n9459
                           , QN => n25272);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n7717, CK => CLK, Q => n9464
                           , QN => n25273);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n7716, CK => CLK, Q => n9469
                           , QN => n25274);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n7715, CK => CLK, Q => n9474
                           , QN => n25275);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n7714, CK => CLK, Q => n9479
                           , QN => n25276);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n7713, CK => CLK, Q => n9484
                           , QN => n25277);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n7712, CK => CLK, Q => n9489
                           , QN => n25278);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n7711, CK => CLK, Q => n9494
                           , QN => n25279);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n7710, CK => CLK, Q => n9499
                           , QN => n25280);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n7709, CK => CLK, Q => n9504
                           , QN => n25281);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n7708, CK => CLK, Q => n9509
                           , QN => n25282);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n7707, CK => CLK, Q => n9514
                           , QN => n25283);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n7706, CK => CLK, Q => n9519
                           , QN => n25284);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n7705, CK => CLK, Q => n9524
                           , QN => n25285);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n7704, CK => CLK, Q => n9529
                           , QN => n25286);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n7703, CK => CLK, Q => n9534
                           , QN => n25287);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n7702, CK => CLK, Q => n9539
                           , QN => n25288);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n7701, CK => CLK, Q => n9544
                           , QN => n25289);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n7700, CK => CLK, Q => n9549
                           , QN => n25290);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n7699, CK => CLK, Q => n9554
                           , QN => n25291);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n7698, CK => CLK, Q => n9559,
                           QN => n25292);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n7697, CK => CLK, Q => n9564,
                           QN => n25293);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n7696, CK => CLK, Q => n9569,
                           QN => n25294);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n7695, CK => CLK, Q => n9574,
                           QN => n25295);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n7694, CK => CLK, Q => n9579,
                           QN => n25296);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n7693, CK => CLK, Q => n9584,
                           QN => n25297);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n7692, CK => CLK, Q => n9589,
                           QN => n25298);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n7691, CK => CLK, Q => n9594,
                           QN => n25299);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n7690, CK => CLK, Q => n9599,
                           QN => n25300);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n7689, CK => CLK, Q => n9604,
                           QN => n25301);
   REGISTERS_reg_13_59_inst : DFF_X1 port map( D => n7044, CK => CLK, Q => 
                           n22238, QN => n25742);
   REGISTERS_reg_13_58_inst : DFF_X1 port map( D => n7043, CK => CLK, Q => 
                           n22237, QN => n25743);
   REGISTERS_reg_13_57_inst : DFF_X1 port map( D => n7042, CK => CLK, Q => 
                           n22236, QN => n25744);
   REGISTERS_reg_13_56_inst : DFF_X1 port map( D => n7041, CK => CLK, Q => 
                           n22235, QN => n25745);
   REGISTERS_reg_13_55_inst : DFF_X1 port map( D => n7040, CK => CLK, Q => 
                           n22234, QN => n25746);
   REGISTERS_reg_13_54_inst : DFF_X1 port map( D => n7039, CK => CLK, Q => 
                           n22233, QN => n25747);
   REGISTERS_reg_13_53_inst : DFF_X1 port map( D => n7038, CK => CLK, Q => 
                           n22232, QN => n25748);
   REGISTERS_reg_13_52_inst : DFF_X1 port map( D => n7037, CK => CLK, Q => 
                           n22231, QN => n25749);
   REGISTERS_reg_13_51_inst : DFF_X1 port map( D => n7036, CK => CLK, Q => 
                           n22230, QN => n25750);
   REGISTERS_reg_13_50_inst : DFF_X1 port map( D => n7035, CK => CLK, Q => 
                           n22229, QN => n25751);
   REGISTERS_reg_13_49_inst : DFF_X1 port map( D => n7034, CK => CLK, Q => 
                           n22228, QN => n25752);
   REGISTERS_reg_13_48_inst : DFF_X1 port map( D => n7033, CK => CLK, Q => 
                           n22227, QN => n25753);
   REGISTERS_reg_13_47_inst : DFF_X1 port map( D => n7032, CK => CLK, Q => 
                           n22226, QN => n25754);
   REGISTERS_reg_13_46_inst : DFF_X1 port map( D => n7031, CK => CLK, Q => 
                           n22225, QN => n25755);
   REGISTERS_reg_13_45_inst : DFF_X1 port map( D => n7030, CK => CLK, Q => 
                           n22224, QN => n25756);
   REGISTERS_reg_13_44_inst : DFF_X1 port map( D => n7029, CK => CLK, Q => 
                           n22223, QN => n25757);
   REGISTERS_reg_13_43_inst : DFF_X1 port map( D => n7028, CK => CLK, Q => 
                           n22222, QN => n25758);
   REGISTERS_reg_13_42_inst : DFF_X1 port map( D => n7027, CK => CLK, Q => 
                           n22221, QN => n25759);
   REGISTERS_reg_13_41_inst : DFF_X1 port map( D => n7026, CK => CLK, Q => 
                           n22220, QN => n25760);
   REGISTERS_reg_13_40_inst : DFF_X1 port map( D => n7025, CK => CLK, Q => 
                           n22219, QN => n25761);
   REGISTERS_reg_13_39_inst : DFF_X1 port map( D => n7024, CK => CLK, Q => 
                           n22218, QN => n25762);
   REGISTERS_reg_13_38_inst : DFF_X1 port map( D => n7023, CK => CLK, Q => 
                           n22217, QN => n25763);
   REGISTERS_reg_13_37_inst : DFF_X1 port map( D => n7022, CK => CLK, Q => 
                           n22216, QN => n25764);
   REGISTERS_reg_13_36_inst : DFF_X1 port map( D => n7021, CK => CLK, Q => 
                           n22215, QN => n25765);
   REGISTERS_reg_13_35_inst : DFF_X1 port map( D => n7020, CK => CLK, Q => 
                           n22214, QN => n25766);
   REGISTERS_reg_13_34_inst : DFF_X1 port map( D => n7019, CK => CLK, Q => 
                           n22213, QN => n25767);
   REGISTERS_reg_13_33_inst : DFF_X1 port map( D => n7018, CK => CLK, Q => 
                           n22212, QN => n25768);
   REGISTERS_reg_13_32_inst : DFF_X1 port map( D => n7017, CK => CLK, Q => 
                           n22211, QN => n25769);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n7016, CK => CLK, Q => 
                           n22210, QN => n25770);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n7015, CK => CLK, Q => 
                           n22209, QN => n25771);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n7014, CK => CLK, Q => 
                           n22208, QN => n25772);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n7013, CK => CLK, Q => 
                           n22207, QN => n25773);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n7012, CK => CLK, Q => 
                           n22206, QN => n25774);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n7011, CK => CLK, Q => 
                           n22205, QN => n25775);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n7010, CK => CLK, Q => 
                           n22204, QN => n25776);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n7009, CK => CLK, Q => 
                           n22203, QN => n25777);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n7008, CK => CLK, Q => 
                           n22202, QN => n25778);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n7007, CK => CLK, Q => 
                           n22201, QN => n25779);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n7006, CK => CLK, Q => 
                           n22200, QN => n25780);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n7005, CK => CLK, Q => 
                           n22199, QN => n25781);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n7004, CK => CLK, Q => 
                           n22198, QN => n25782);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n7003, CK => CLK, Q => 
                           n22197, QN => n25783);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n7002, CK => CLK, Q => 
                           n22196, QN => n25784);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n7001, CK => CLK, Q => 
                           n22195, QN => n25785);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n7000, CK => CLK, Q => 
                           n22194, QN => n25786);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n6999, CK => CLK, Q => 
                           n22193, QN => n25787);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n6998, CK => CLK, Q => 
                           n22192, QN => n25788);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n6997, CK => CLK, Q => 
                           n22191, QN => n25789);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n6996, CK => CLK, Q => 
                           n22190, QN => n25790);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n6995, CK => CLK, Q => 
                           n22189, QN => n25791);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n6994, CK => CLK, Q => 
                           n22188, QN => n25792);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n6993, CK => CLK, Q => 
                           n22187, QN => n25793);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n6992, CK => CLK, Q => 
                           n22186, QN => n25794);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n6991, CK => CLK, Q => 
                           n22185, QN => n25795);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n6990, CK => CLK, Q => 
                           n22184, QN => n25796);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n6989, CK => CLK, Q => 
                           n22183, QN => n25797);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n6988, CK => CLK, Q => 
                           n22182, QN => n25798);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n6987, CK => CLK, Q => 
                           n22181, QN => n25799);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n6986, CK => CLK, Q => 
                           n22180, QN => n25800);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n6985, CK => CLK, Q => 
                           n22179, QN => n25801);
   REGISTERS_reg_9_59_inst : DFF_X1 port map( D => n7300, CK => CLK, Q => 
                           n21986, QN => n25594);
   REGISTERS_reg_9_58_inst : DFF_X1 port map( D => n7299, CK => CLK, Q => 
                           n21985, QN => n25595);
   REGISTERS_reg_9_57_inst : DFF_X1 port map( D => n7298, CK => CLK, Q => 
                           n21984, QN => n25596);
   REGISTERS_reg_9_56_inst : DFF_X1 port map( D => n7297, CK => CLK, Q => 
                           n21983, QN => n25597);
   REGISTERS_reg_9_55_inst : DFF_X1 port map( D => n7296, CK => CLK, Q => 
                           n21982, QN => n25598);
   REGISTERS_reg_9_54_inst : DFF_X1 port map( D => n7295, CK => CLK, Q => 
                           n21981, QN => n25599);
   REGISTERS_reg_9_53_inst : DFF_X1 port map( D => n7294, CK => CLK, Q => 
                           n21980, QN => n25600);
   REGISTERS_reg_9_52_inst : DFF_X1 port map( D => n7293, CK => CLK, Q => 
                           n21979, QN => n25601);
   REGISTERS_reg_9_51_inst : DFF_X1 port map( D => n7292, CK => CLK, Q => 
                           n21978, QN => n25602);
   REGISTERS_reg_9_50_inst : DFF_X1 port map( D => n7291, CK => CLK, Q => 
                           n21977, QN => n25603);
   REGISTERS_reg_9_49_inst : DFF_X1 port map( D => n7290, CK => CLK, Q => 
                           n21976, QN => n25604);
   REGISTERS_reg_9_48_inst : DFF_X1 port map( D => n7289, CK => CLK, Q => 
                           n21975, QN => n25605);
   REGISTERS_reg_9_47_inst : DFF_X1 port map( D => n7288, CK => CLK, Q => 
                           n21974, QN => n25606);
   REGISTERS_reg_9_46_inst : DFF_X1 port map( D => n7287, CK => CLK, Q => 
                           n21973, QN => n25607);
   REGISTERS_reg_9_45_inst : DFF_X1 port map( D => n7286, CK => CLK, Q => 
                           n21972, QN => n25608);
   REGISTERS_reg_9_44_inst : DFF_X1 port map( D => n7285, CK => CLK, Q => 
                           n21971, QN => n25609);
   REGISTERS_reg_9_43_inst : DFF_X1 port map( D => n7284, CK => CLK, Q => 
                           n21970, QN => n25610);
   REGISTERS_reg_9_42_inst : DFF_X1 port map( D => n7283, CK => CLK, Q => 
                           n21969, QN => n25611);
   REGISTERS_reg_9_41_inst : DFF_X1 port map( D => n7282, CK => CLK, Q => 
                           n21968, QN => n25612);
   REGISTERS_reg_9_40_inst : DFF_X1 port map( D => n7281, CK => CLK, Q => 
                           n21967, QN => n25613);
   REGISTERS_reg_9_39_inst : DFF_X1 port map( D => n7280, CK => CLK, Q => 
                           n21966, QN => n25614);
   REGISTERS_reg_9_38_inst : DFF_X1 port map( D => n7279, CK => CLK, Q => 
                           n21965, QN => n25615);
   REGISTERS_reg_9_37_inst : DFF_X1 port map( D => n7278, CK => CLK, Q => 
                           n21964, QN => n25616);
   REGISTERS_reg_9_36_inst : DFF_X1 port map( D => n7277, CK => CLK, Q => 
                           n21963, QN => n25617);
   REGISTERS_reg_9_35_inst : DFF_X1 port map( D => n7276, CK => CLK, Q => 
                           n21962, QN => n25618);
   REGISTERS_reg_9_34_inst : DFF_X1 port map( D => n7275, CK => CLK, Q => 
                           n21961, QN => n25619);
   REGISTERS_reg_9_33_inst : DFF_X1 port map( D => n7274, CK => CLK, Q => 
                           n21960, QN => n25620);
   REGISTERS_reg_9_32_inst : DFF_X1 port map( D => n7273, CK => CLK, Q => 
                           n21959, QN => n25621);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n7272, CK => CLK, Q => 
                           n21958, QN => n25622);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n7271, CK => CLK, Q => 
                           n21957, QN => n25623);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n7270, CK => CLK, Q => 
                           n21956, QN => n25624);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n7269, CK => CLK, Q => 
                           n21955, QN => n25625);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n7268, CK => CLK, Q => 
                           n21954, QN => n25626);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n7267, CK => CLK, Q => 
                           n21953, QN => n25627);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n7266, CK => CLK, Q => 
                           n21952, QN => n25628);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n7265, CK => CLK, Q => 
                           n21951, QN => n25629);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n7264, CK => CLK, Q => 
                           n21950, QN => n25630);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n7263, CK => CLK, Q => 
                           n21949, QN => n25631);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n7262, CK => CLK, Q => 
                           n21948, QN => n25632);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n7261, CK => CLK, Q => 
                           n21947, QN => n25633);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n7260, CK => CLK, Q => 
                           n21946, QN => n25634);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n7259, CK => CLK, Q => 
                           n21945, QN => n25635);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n7258, CK => CLK, Q => 
                           n21944, QN => n25636);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n7257, CK => CLK, Q => 
                           n21943, QN => n25637);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n7256, CK => CLK, Q => 
                           n21942, QN => n25638);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n7255, CK => CLK, Q => 
                           n21941, QN => n25639);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n7254, CK => CLK, Q => 
                           n21940, QN => n25640);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n7253, CK => CLK, Q => 
                           n21939, QN => n25641);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n7252, CK => CLK, Q => 
                           n21938, QN => n25642);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n7251, CK => CLK, Q => 
                           n21937, QN => n25643);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n7250, CK => CLK, Q => n21936
                           , QN => n25644);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n7249, CK => CLK, Q => n21935
                           , QN => n25645);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n7248, CK => CLK, Q => n21934
                           , QN => n25646);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n7247, CK => CLK, Q => n21933
                           , QN => n25647);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n7246, CK => CLK, Q => n21932
                           , QN => n25648);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n7245, CK => CLK, Q => n21931
                           , QN => n25649);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n7244, CK => CLK, Q => n21930
                           , QN => n25650);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n7243, CK => CLK, Q => n21929
                           , QN => n25651);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n7242, CK => CLK, Q => n21928
                           , QN => n25652);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n7241, CK => CLK, Q => n21927
                           , QN => n25653);
   REGISTERS_reg_7_59_inst : DFF_X1 port map( D => n7428, CK => CLK, Q => 
                           n22064, QN => n25461);
   REGISTERS_reg_7_58_inst : DFF_X1 port map( D => n7427, CK => CLK, Q => 
                           n22063, QN => n25462);
   REGISTERS_reg_7_57_inst : DFF_X1 port map( D => n7426, CK => CLK, Q => 
                           n22062, QN => n25463);
   REGISTERS_reg_7_56_inst : DFF_X1 port map( D => n7425, CK => CLK, Q => 
                           n22061, QN => n25464);
   REGISTERS_reg_7_55_inst : DFF_X1 port map( D => n7424, CK => CLK, Q => 
                           n22060, QN => n25465);
   REGISTERS_reg_7_54_inst : DFF_X1 port map( D => n7423, CK => CLK, Q => 
                           n22059, QN => n25466);
   REGISTERS_reg_7_53_inst : DFF_X1 port map( D => n7422, CK => CLK, Q => 
                           n22058, QN => n25467);
   REGISTERS_reg_7_52_inst : DFF_X1 port map( D => n7421, CK => CLK, Q => 
                           n22057, QN => n25468);
   REGISTERS_reg_7_51_inst : DFF_X1 port map( D => n7420, CK => CLK, Q => 
                           n22056, QN => n25469);
   REGISTERS_reg_7_50_inst : DFF_X1 port map( D => n7419, CK => CLK, Q => 
                           n22055, QN => n25470);
   REGISTERS_reg_7_49_inst : DFF_X1 port map( D => n7418, CK => CLK, Q => 
                           n22054, QN => n25471);
   REGISTERS_reg_7_48_inst : DFF_X1 port map( D => n7417, CK => CLK, Q => 
                           n22053, QN => n25472);
   REGISTERS_reg_7_47_inst : DFF_X1 port map( D => n7416, CK => CLK, Q => 
                           n22052, QN => n25473);
   REGISTERS_reg_7_46_inst : DFF_X1 port map( D => n7415, CK => CLK, Q => 
                           n22051, QN => n25474);
   REGISTERS_reg_7_45_inst : DFF_X1 port map( D => n7414, CK => CLK, Q => 
                           n22050, QN => n25475);
   REGISTERS_reg_7_44_inst : DFF_X1 port map( D => n7413, CK => CLK, Q => 
                           n22049, QN => n25476);
   REGISTERS_reg_7_43_inst : DFF_X1 port map( D => n7412, CK => CLK, Q => 
                           n22048, QN => n25477);
   REGISTERS_reg_7_42_inst : DFF_X1 port map( D => n7411, CK => CLK, Q => 
                           n22047, QN => n25478);
   REGISTERS_reg_7_41_inst : DFF_X1 port map( D => n7410, CK => CLK, Q => 
                           n22046, QN => n25479);
   REGISTERS_reg_7_40_inst : DFF_X1 port map( D => n7409, CK => CLK, Q => 
                           n22045, QN => n25480);
   REGISTERS_reg_7_39_inst : DFF_X1 port map( D => n7408, CK => CLK, Q => 
                           n22044, QN => n25481);
   REGISTERS_reg_7_38_inst : DFF_X1 port map( D => n7407, CK => CLK, Q => 
                           n22043, QN => n25482);
   REGISTERS_reg_7_37_inst : DFF_X1 port map( D => n7406, CK => CLK, Q => 
                           n22042, QN => n25483);
   REGISTERS_reg_7_36_inst : DFF_X1 port map( D => n7405, CK => CLK, Q => 
                           n22041, QN => n25484);
   REGISTERS_reg_7_35_inst : DFF_X1 port map( D => n7404, CK => CLK, Q => 
                           n22040, QN => n25485);
   REGISTERS_reg_7_34_inst : DFF_X1 port map( D => n7403, CK => CLK, Q => 
                           n22039, QN => n25486);
   REGISTERS_reg_7_33_inst : DFF_X1 port map( D => n7402, CK => CLK, Q => 
                           n22038, QN => n25487);
   REGISTERS_reg_7_32_inst : DFF_X1 port map( D => n7401, CK => CLK, Q => 
                           n22037, QN => n25488);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n7400, CK => CLK, Q => 
                           n22036, QN => n25489);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n7399, CK => CLK, Q => 
                           n22035, QN => n25490);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n7398, CK => CLK, Q => 
                           n22034, QN => n25491);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n7397, CK => CLK, Q => 
                           n22033, QN => n25492);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n7396, CK => CLK, Q => 
                           n22032, QN => n25493);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n7395, CK => CLK, Q => 
                           n22031, QN => n25494);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n7394, CK => CLK, Q => 
                           n22030, QN => n25495);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n7393, CK => CLK, Q => 
                           n22029, QN => n25496);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n7392, CK => CLK, Q => 
                           n22028, QN => n25497);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n7391, CK => CLK, Q => 
                           n22027, QN => n25498);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n7390, CK => CLK, Q => 
                           n22026, QN => n25499);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n7389, CK => CLK, Q => 
                           n22025, QN => n25500);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n7388, CK => CLK, Q => 
                           n22024, QN => n25501);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n7387, CK => CLK, Q => 
                           n22023, QN => n25502);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n7386, CK => CLK, Q => 
                           n22022, QN => n25503);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n7385, CK => CLK, Q => 
                           n22021, QN => n25504);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n7384, CK => CLK, Q => 
                           n22020, QN => n25505);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n7383, CK => CLK, Q => 
                           n22019, QN => n25506);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n7382, CK => CLK, Q => 
                           n22018, QN => n25507);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n7381, CK => CLK, Q => 
                           n22017, QN => n25508);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n7380, CK => CLK, Q => 
                           n22016, QN => n25509);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n7379, CK => CLK, Q => 
                           n22075, QN => n25510);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n7378, CK => CLK, Q => n22074
                           , QN => n25511);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n7377, CK => CLK, Q => n22073
                           , QN => n25512);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n7376, CK => CLK, Q => n22072
                           , QN => n25513);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n7375, CK => CLK, Q => n22071
                           , QN => n25514);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n7374, CK => CLK, Q => n22070
                           , QN => n25515);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n7373, CK => CLK, Q => n22069
                           , QN => n25516);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n7372, CK => CLK, Q => n22068
                           , QN => n25517);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n7371, CK => CLK, Q => n22067
                           , QN => n25518);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n7370, CK => CLK, Q => n22066
                           , QN => n25519);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n7369, CK => CLK, Q => n22065
                           , QN => n25520);
   REGISTERS_reg_3_59_inst : DFF_X1 port map( D => n7684, CK => CLK, Q => 
                           n21854, QN => n25309);
   REGISTERS_reg_3_58_inst : DFF_X1 port map( D => n7683, CK => CLK, Q => 
                           n21853, QN => n25310);
   REGISTERS_reg_3_57_inst : DFF_X1 port map( D => n7682, CK => CLK, Q => 
                           n21852, QN => n25311);
   REGISTERS_reg_3_56_inst : DFF_X1 port map( D => n7681, CK => CLK, Q => 
                           n21851, QN => n25312);
   REGISTERS_reg_3_55_inst : DFF_X1 port map( D => n7680, CK => CLK, Q => 
                           n21850, QN => n25313);
   REGISTERS_reg_3_54_inst : DFF_X1 port map( D => n7679, CK => CLK, Q => 
                           n21849, QN => n25314);
   REGISTERS_reg_3_53_inst : DFF_X1 port map( D => n7678, CK => CLK, Q => 
                           n21848, QN => n25315);
   REGISTERS_reg_3_52_inst : DFF_X1 port map( D => n7677, CK => CLK, Q => 
                           n21847, QN => n25316);
   REGISTERS_reg_3_51_inst : DFF_X1 port map( D => n7676, CK => CLK, Q => 
                           n21846, QN => n25317);
   REGISTERS_reg_3_50_inst : DFF_X1 port map( D => n7675, CK => CLK, Q => 
                           n21845, QN => n25318);
   REGISTERS_reg_3_49_inst : DFF_X1 port map( D => n7674, CK => CLK, Q => 
                           n21844, QN => n25319);
   REGISTERS_reg_3_48_inst : DFF_X1 port map( D => n7673, CK => CLK, Q => 
                           n21843, QN => n25320);
   REGISTERS_reg_3_47_inst : DFF_X1 port map( D => n7672, CK => CLK, Q => 
                           n21842, QN => n25321);
   REGISTERS_reg_3_46_inst : DFF_X1 port map( D => n7671, CK => CLK, Q => 
                           n21841, QN => n25322);
   REGISTERS_reg_3_45_inst : DFF_X1 port map( D => n7670, CK => CLK, Q => 
                           n21840, QN => n25323);
   REGISTERS_reg_3_44_inst : DFF_X1 port map( D => n7669, CK => CLK, Q => 
                           n21839, QN => n25324);
   REGISTERS_reg_3_43_inst : DFF_X1 port map( D => n7668, CK => CLK, Q => 
                           n21838, QN => n25325);
   REGISTERS_reg_3_42_inst : DFF_X1 port map( D => n7667, CK => CLK, Q => 
                           n21837, QN => n25326);
   REGISTERS_reg_3_41_inst : DFF_X1 port map( D => n7666, CK => CLK, Q => 
                           n21836, QN => n25327);
   REGISTERS_reg_3_40_inst : DFF_X1 port map( D => n7665, CK => CLK, Q => 
                           n21835, QN => n25328);
   REGISTERS_reg_3_39_inst : DFF_X1 port map( D => n7664, CK => CLK, Q => 
                           n21834, QN => n25329);
   REGISTERS_reg_3_38_inst : DFF_X1 port map( D => n7663, CK => CLK, Q => 
                           n21833, QN => n25330);
   REGISTERS_reg_3_37_inst : DFF_X1 port map( D => n7662, CK => CLK, Q => 
                           n21832, QN => n25331);
   REGISTERS_reg_3_36_inst : DFF_X1 port map( D => n7661, CK => CLK, Q => 
                           n21831, QN => n25332);
   REGISTERS_reg_3_35_inst : DFF_X1 port map( D => n7660, CK => CLK, Q => 
                           n21830, QN => n25333);
   REGISTERS_reg_3_34_inst : DFF_X1 port map( D => n7659, CK => CLK, Q => 
                           n21829, QN => n25334);
   REGISTERS_reg_3_33_inst : DFF_X1 port map( D => n7658, CK => CLK, Q => 
                           n21828, QN => n25335);
   REGISTERS_reg_3_32_inst : DFF_X1 port map( D => n7657, CK => CLK, Q => 
                           n21827, QN => n25336);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n7656, CK => CLK, Q => 
                           n21826, QN => n25337);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n7655, CK => CLK, Q => 
                           n21825, QN => n25338);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n7654, CK => CLK, Q => 
                           n21824, QN => n25339);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n7653, CK => CLK, Q => 
                           n21823, QN => n25340);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n7652, CK => CLK, Q => 
                           n21822, QN => n25341);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n7651, CK => CLK, Q => 
                           n21821, QN => n25342);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n7650, CK => CLK, Q => 
                           n21820, QN => n25343);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n7649, CK => CLK, Q => 
                           n21819, QN => n25344);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n7648, CK => CLK, Q => 
                           n21818, QN => n25345);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n7647, CK => CLK, Q => 
                           n21817, QN => n25346);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n7646, CK => CLK, Q => 
                           n21816, QN => n25347);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n7645, CK => CLK, Q => 
                           n21815, QN => n25348);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n7644, CK => CLK, Q => 
                           n21814, QN => n25349);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n7643, CK => CLK, Q => 
                           n21813, QN => n25350);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n7642, CK => CLK, Q => 
                           n21812, QN => n25351);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n7641, CK => CLK, Q => 
                           n21811, QN => n25352);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n7640, CK => CLK, Q => 
                           n21810, QN => n25353);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n7639, CK => CLK, Q => 
                           n21809, QN => n25354);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n7638, CK => CLK, Q => 
                           n21808, QN => n25355);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n7637, CK => CLK, Q => 
                           n21807, QN => n25356);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n7636, CK => CLK, Q => 
                           n21806, QN => n25357);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n7635, CK => CLK, Q => 
                           n21805, QN => n25358);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n7634, CK => CLK, Q => n21804
                           , QN => n25359);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n7633, CK => CLK, Q => n21803
                           , QN => n25360);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n7632, CK => CLK, Q => n21802
                           , QN => n25361);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n7631, CK => CLK, Q => n21801
                           , QN => n25362);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n7630, CK => CLK, Q => n21800
                           , QN => n25363);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n7629, CK => CLK, Q => n21799
                           , QN => n25364);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n7628, CK => CLK, Q => n21798
                           , QN => n25365);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n7627, CK => CLK, Q => n21797
                           , QN => n25366);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n7626, CK => CLK, Q => n21796
                           , QN => n25367);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n7625, CK => CLK, Q => n21795
                           , QN => n25368);
   REGISTERS_reg_12_59_inst : DFF_X1 port map( D => n7108, CK => CLK, Q => 
                           n9677, QN => n25676);
   REGISTERS_reg_12_58_inst : DFF_X1 port map( D => n7107, CK => CLK, Q => 
                           n9678, QN => n25677);
   REGISTERS_reg_12_57_inst : DFF_X1 port map( D => n7106, CK => CLK, Q => 
                           n9679, QN => n25678);
   REGISTERS_reg_12_56_inst : DFF_X1 port map( D => n7105, CK => CLK, Q => 
                           n9680, QN => n25679);
   REGISTERS_reg_12_55_inst : DFF_X1 port map( D => n7104, CK => CLK, Q => 
                           n9681, QN => n25680);
   REGISTERS_reg_12_54_inst : DFF_X1 port map( D => n7103, CK => CLK, Q => 
                           n9682, QN => n25681);
   REGISTERS_reg_12_53_inst : DFF_X1 port map( D => n7102, CK => CLK, Q => 
                           n9683, QN => n25682);
   REGISTERS_reg_12_52_inst : DFF_X1 port map( D => n7101, CK => CLK, Q => 
                           n9684, QN => n25683);
   REGISTERS_reg_12_51_inst : DFF_X1 port map( D => n7100, CK => CLK, Q => 
                           n9685, QN => n25684);
   REGISTERS_reg_12_50_inst : DFF_X1 port map( D => n7099, CK => CLK, Q => 
                           n9686, QN => n25685);
   REGISTERS_reg_12_49_inst : DFF_X1 port map( D => n7098, CK => CLK, Q => 
                           n9687, QN => n25686);
   REGISTERS_reg_12_48_inst : DFF_X1 port map( D => n7097, CK => CLK, Q => 
                           n9688, QN => n25687);
   REGISTERS_reg_12_47_inst : DFF_X1 port map( D => n7096, CK => CLK, Q => 
                           n9689, QN => n25688);
   REGISTERS_reg_12_46_inst : DFF_X1 port map( D => n7095, CK => CLK, Q => 
                           n9690, QN => n25689);
   REGISTERS_reg_12_45_inst : DFF_X1 port map( D => n7094, CK => CLK, Q => 
                           n9691, QN => n25690);
   REGISTERS_reg_12_44_inst : DFF_X1 port map( D => n7093, CK => CLK, Q => 
                           n9692, QN => n25691);
   REGISTERS_reg_12_43_inst : DFF_X1 port map( D => n7092, CK => CLK, Q => 
                           n9693, QN => n25692);
   REGISTERS_reg_12_42_inst : DFF_X1 port map( D => n7091, CK => CLK, Q => 
                           n9694, QN => n25693);
   REGISTERS_reg_12_41_inst : DFF_X1 port map( D => n7090, CK => CLK, Q => 
                           n9695, QN => n25694);
   REGISTERS_reg_12_40_inst : DFF_X1 port map( D => n7089, CK => CLK, Q => 
                           n9696, QN => n25695);
   REGISTERS_reg_12_39_inst : DFF_X1 port map( D => n7088, CK => CLK, Q => 
                           n9697, QN => n25696);
   REGISTERS_reg_12_38_inst : DFF_X1 port map( D => n7087, CK => CLK, Q => 
                           n9698, QN => n25697);
   REGISTERS_reg_12_37_inst : DFF_X1 port map( D => n7086, CK => CLK, Q => 
                           n9699, QN => n25698);
   REGISTERS_reg_12_36_inst : DFF_X1 port map( D => n7085, CK => CLK, Q => 
                           n9700, QN => n25699);
   REGISTERS_reg_12_35_inst : DFF_X1 port map( D => n7084, CK => CLK, Q => 
                           n9701, QN => n25700);
   REGISTERS_reg_12_34_inst : DFF_X1 port map( D => n7083, CK => CLK, Q => 
                           n9702, QN => n25701);
   REGISTERS_reg_12_33_inst : DFF_X1 port map( D => n7082, CK => CLK, Q => 
                           n9703, QN => n25702);
   REGISTERS_reg_12_32_inst : DFF_X1 port map( D => n7081, CK => CLK, Q => 
                           n9704, QN => n25703);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n7080, CK => CLK, Q => 
                           n9705, QN => n25704);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n7079, CK => CLK, Q => 
                           n9706, QN => n25705);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n7078, CK => CLK, Q => 
                           n9707, QN => n25706);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n7077, CK => CLK, Q => 
                           n9708, QN => n25707);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n7076, CK => CLK, Q => 
                           n9709, QN => n25708);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n7075, CK => CLK, Q => 
                           n9710, QN => n25709);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n7074, CK => CLK, Q => 
                           n9711, QN => n25710);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n7073, CK => CLK, Q => 
                           n9712, QN => n25711);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n7072, CK => CLK, Q => 
                           n9713, QN => n25712);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n7071, CK => CLK, Q => 
                           n9714, QN => n25713);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n7070, CK => CLK, Q => 
                           n9715, QN => n25714);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n7069, CK => CLK, Q => 
                           n9716, QN => n25715);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n7068, CK => CLK, Q => 
                           n9717, QN => n25716);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n7067, CK => CLK, Q => 
                           n9718, QN => n25717);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n7066, CK => CLK, Q => 
                           n9719, QN => n25718);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n7065, CK => CLK, Q => 
                           n9720, QN => n25719);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n7064, CK => CLK, Q => 
                           n9721, QN => n25720);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n7063, CK => CLK, Q => 
                           n9722, QN => n25721);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n7062, CK => CLK, Q => 
                           n9723, QN => n25722);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n7061, CK => CLK, Q => 
                           n9724, QN => n25723);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n7060, CK => CLK, Q => 
                           n9725, QN => n25724);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n7059, CK => CLK, Q => 
                           n9726, QN => n25725);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n7058, CK => CLK, Q => n9727
                           , QN => n25726);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n7057, CK => CLK, Q => n9728
                           , QN => n25727);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n7056, CK => CLK, Q => n9729
                           , QN => n25728);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n7055, CK => CLK, Q => n9730
                           , QN => n25729);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n7054, CK => CLK, Q => n9731
                           , QN => n25730);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n7053, CK => CLK, Q => n9732
                           , QN => n25731);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n7052, CK => CLK, Q => n9733
                           , QN => n25732);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n7051, CK => CLK, Q => n9734
                           , QN => n25733);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n7050, CK => CLK, Q => n9735
                           , QN => n25734);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n7049, CK => CLK, Q => n9736
                           , QN => n25735);
   REGISTERS_reg_8_59_inst : DFF_X1 port map( D => n7364, CK => CLK, Q => n9311
                           , QN => n25527);
   REGISTERS_reg_8_58_inst : DFF_X1 port map( D => n7363, CK => CLK, Q => n9316
                           , QN => n25528);
   REGISTERS_reg_8_57_inst : DFF_X1 port map( D => n7362, CK => CLK, Q => n9321
                           , QN => n25529);
   REGISTERS_reg_8_56_inst : DFF_X1 port map( D => n7361, CK => CLK, Q => n9326
                           , QN => n25530);
   REGISTERS_reg_8_55_inst : DFF_X1 port map( D => n7360, CK => CLK, Q => n9331
                           , QN => n25531);
   REGISTERS_reg_8_54_inst : DFF_X1 port map( D => n7359, CK => CLK, Q => n9336
                           , QN => n25532);
   REGISTERS_reg_8_53_inst : DFF_X1 port map( D => n7358, CK => CLK, Q => n9341
                           , QN => n25533);
   REGISTERS_reg_8_52_inst : DFF_X1 port map( D => n7357, CK => CLK, Q => n9346
                           , QN => n25534);
   REGISTERS_reg_8_51_inst : DFF_X1 port map( D => n7356, CK => CLK, Q => n9351
                           , QN => n25535);
   REGISTERS_reg_8_50_inst : DFF_X1 port map( D => n7355, CK => CLK, Q => n9356
                           , QN => n25536);
   REGISTERS_reg_8_49_inst : DFF_X1 port map( D => n7354, CK => CLK, Q => n9361
                           , QN => n25537);
   REGISTERS_reg_8_48_inst : DFF_X1 port map( D => n7353, CK => CLK, Q => n9366
                           , QN => n25538);
   REGISTERS_reg_8_47_inst : DFF_X1 port map( D => n7352, CK => CLK, Q => n9371
                           , QN => n25539);
   REGISTERS_reg_8_46_inst : DFF_X1 port map( D => n7351, CK => CLK, Q => n9376
                           , QN => n25540);
   REGISTERS_reg_8_45_inst : DFF_X1 port map( D => n7350, CK => CLK, Q => n9381
                           , QN => n25541);
   REGISTERS_reg_8_44_inst : DFF_X1 port map( D => n7349, CK => CLK, Q => n9386
                           , QN => n25542);
   REGISTERS_reg_8_43_inst : DFF_X1 port map( D => n7348, CK => CLK, Q => n9391
                           , QN => n25543);
   REGISTERS_reg_8_42_inst : DFF_X1 port map( D => n7347, CK => CLK, Q => n9396
                           , QN => n25544);
   REGISTERS_reg_8_41_inst : DFF_X1 port map( D => n7346, CK => CLK, Q => n9401
                           , QN => n25545);
   REGISTERS_reg_8_40_inst : DFF_X1 port map( D => n7345, CK => CLK, Q => n9406
                           , QN => n25546);
   REGISTERS_reg_8_39_inst : DFF_X1 port map( D => n7344, CK => CLK, Q => n9411
                           , QN => n25547);
   REGISTERS_reg_8_38_inst : DFF_X1 port map( D => n7343, CK => CLK, Q => n9416
                           , QN => n25548);
   REGISTERS_reg_8_37_inst : DFF_X1 port map( D => n7342, CK => CLK, Q => n9421
                           , QN => n25549);
   REGISTERS_reg_8_36_inst : DFF_X1 port map( D => n7341, CK => CLK, Q => n9426
                           , QN => n25550);
   REGISTERS_reg_8_35_inst : DFF_X1 port map( D => n7340, CK => CLK, Q => n9431
                           , QN => n25551);
   REGISTERS_reg_8_34_inst : DFF_X1 port map( D => n7339, CK => CLK, Q => n9436
                           , QN => n25552);
   REGISTERS_reg_8_33_inst : DFF_X1 port map( D => n7338, CK => CLK, Q => n9441
                           , QN => n25553);
   REGISTERS_reg_8_32_inst : DFF_X1 port map( D => n7337, CK => CLK, Q => n9446
                           , QN => n25554);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n7336, CK => CLK, Q => n9451
                           , QN => n25555);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n7335, CK => CLK, Q => n9456
                           , QN => n25556);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n7334, CK => CLK, Q => n9461
                           , QN => n25557);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n7333, CK => CLK, Q => n9466
                           , QN => n25558);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n7332, CK => CLK, Q => n9471
                           , QN => n25559);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n7331, CK => CLK, Q => n9476
                           , QN => n25560);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n7330, CK => CLK, Q => n9481
                           , QN => n25561);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n7329, CK => CLK, Q => n9486
                           , QN => n25562);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n7328, CK => CLK, Q => n9491
                           , QN => n25563);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n7327, CK => CLK, Q => n9496
                           , QN => n25564);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n7326, CK => CLK, Q => n9501
                           , QN => n25565);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n7325, CK => CLK, Q => n9506
                           , QN => n25566);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n7324, CK => CLK, Q => n9511
                           , QN => n25567);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n7323, CK => CLK, Q => n9516
                           , QN => n25568);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n7322, CK => CLK, Q => n9521
                           , QN => n25569);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n7321, CK => CLK, Q => n9526
                           , QN => n25570);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n7320, CK => CLK, Q => n9531
                           , QN => n25571);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n7319, CK => CLK, Q => n9536
                           , QN => n25572);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n7318, CK => CLK, Q => n9541
                           , QN => n25573);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n7317, CK => CLK, Q => n9546
                           , QN => n25574);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n7316, CK => CLK, Q => n9551
                           , QN => n25575);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n7315, CK => CLK, Q => n9556
                           , QN => n25576);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n7314, CK => CLK, Q => n9561,
                           QN => n25577);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n7313, CK => CLK, Q => n9566,
                           QN => n25578);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n7312, CK => CLK, Q => n9571,
                           QN => n25579);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n7311, CK => CLK, Q => n9576,
                           QN => n25580);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n7310, CK => CLK, Q => n9581,
                           QN => n25581);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n7309, CK => CLK, Q => n9586,
                           QN => n25582);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n7308, CK => CLK, Q => n9591,
                           QN => n25583);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n7307, CK => CLK, Q => n9596,
                           QN => n25584);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n7306, CK => CLK, Q => n9601,
                           QN => n25585);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n7305, CK => CLK, Q => n9606,
                           QN => n25586);
   U19730 : NOR2_X1 port map( A1 => n29305, A2 => ADD_RD1(1), ZN => n29286);
   U19731 : NOR2_X1 port map( A1 => n28028, A2 => ADD_RD2(1), ZN => n28005);
   U19732 : BUF_X1 port map( A => n25155, Z => n31137);
   U19733 : BUF_X1 port map( A => n25155, Z => n31138);
   U19734 : BUF_X1 port map( A => n25155, Z => n31139);
   U19735 : BUF_X1 port map( A => n25155, Z => n31140);
   U19736 : BUF_X1 port map( A => n25523, Z => n30843);
   U19737 : BUF_X1 port map( A => n25523, Z => n30844);
   U19738 : BUF_X1 port map( A => n25523, Z => n30845);
   U19739 : BUF_X1 port map( A => n25523, Z => n30846);
   U19740 : BUF_X1 port map( A => n25523, Z => n30847);
   U19741 : BUF_X1 port map( A => n25672, Z => n30793);
   U19742 : BUF_X1 port map( A => n25672, Z => n30794);
   U19743 : BUF_X1 port map( A => n25672, Z => n30795);
   U19744 : BUF_X1 port map( A => n25672, Z => n30796);
   U19745 : BUF_X1 port map( A => n25672, Z => n30797);
   U19746 : BUF_X1 port map( A => n25238, Z => n30919);
   U19747 : BUF_X1 port map( A => n25238, Z => n30920);
   U19748 : BUF_X1 port map( A => n25238, Z => n30921);
   U19749 : BUF_X1 port map( A => n25238, Z => n30922);
   U19750 : BUF_X1 port map( A => n25238, Z => n30923);
   U19751 : BUF_X1 port map( A => n25387, Z => n30869);
   U19752 : BUF_X1 port map( A => n25387, Z => n30870);
   U19753 : BUF_X1 port map( A => n25387, Z => n30871);
   U19754 : BUF_X1 port map( A => n25387, Z => n30872);
   U19755 : BUF_X1 port map( A => n25387, Z => n30873);
   U19756 : BUF_X1 port map( A => n25809, Z => n30744);
   U19757 : BUF_X1 port map( A => n25809, Z => n30745);
   U19758 : BUF_X1 port map( A => n25809, Z => n30746);
   U19759 : BUF_X1 port map( A => n25809, Z => n30747);
   U19760 : BUF_X1 port map( A => n25809, Z => n30743);
   U19761 : BUF_X1 port map( A => n25959, Z => n30694);
   U19762 : BUF_X1 port map( A => n25959, Z => n30695);
   U19763 : BUF_X1 port map( A => n26025, Z => n30681);
   U19764 : BUF_X1 port map( A => n26025, Z => n30682);
   U19765 : BUF_X1 port map( A => n26104, Z => n30620);
   U19766 : BUF_X1 port map( A => n26104, Z => n30621);
   U19767 : BUF_X1 port map( A => n25959, Z => n30696);
   U19768 : BUF_X1 port map( A => n25959, Z => n30697);
   U19769 : BUF_X1 port map( A => n26025, Z => n30683);
   U19770 : BUF_X1 port map( A => n26025, Z => n30684);
   U19771 : BUF_X1 port map( A => n26104, Z => n30622);
   U19772 : BUF_X1 port map( A => n26104, Z => n30623);
   U19773 : BUF_X1 port map( A => n26252, Z => n30570);
   U19774 : BUF_X1 port map( A => n26252, Z => n30571);
   U19775 : BUF_X1 port map( A => n26252, Z => n30572);
   U19776 : BUF_X1 port map( A => n26252, Z => n30573);
   U19777 : BUF_X1 port map( A => n26318, Z => n30557);
   U19778 : BUF_X1 port map( A => n26318, Z => n30558);
   U19779 : BUF_X1 port map( A => n26318, Z => n30559);
   U19780 : BUF_X1 port map( A => n26318, Z => n30560);
   U19781 : BUF_X1 port map( A => n25959, Z => n30693);
   U19782 : BUF_X1 port map( A => n26025, Z => n30680);
   U19783 : BUF_X1 port map( A => n26104, Z => n30619);
   U19784 : BUF_X1 port map( A => n26252, Z => n30569);
   U19785 : BUF_X1 port map( A => n26318, Z => n30556);
   U19786 : BUF_X1 port map( A => n26170, Z => n30606);
   U19787 : BUF_X1 port map( A => n26170, Z => n30607);
   U19788 : BUF_X1 port map( A => n26170, Z => n30608);
   U19789 : BUF_X1 port map( A => n26170, Z => n30609);
   U19790 : BUF_X1 port map( A => n26170, Z => n30610);
   U19791 : BUF_X1 port map( A => n25876, Z => n30730);
   U19792 : BUF_X1 port map( A => n25876, Z => n30731);
   U19793 : BUF_X1 port map( A => n25876, Z => n30732);
   U19794 : BUF_X1 port map( A => n25876, Z => n30733);
   U19795 : BUF_X1 port map( A => n25876, Z => n30734);
   U19796 : BUF_X1 port map( A => n25738, Z => n30780);
   U19797 : BUF_X1 port map( A => n25738, Z => n30781);
   U19798 : BUF_X1 port map( A => n25738, Z => n30782);
   U19799 : BUF_X1 port map( A => n25738, Z => n30783);
   U19800 : BUF_X1 port map( A => n25738, Z => n30784);
   U19801 : BUF_X1 port map( A => n25590, Z => n30830);
   U19802 : BUF_X1 port map( A => n25590, Z => n30831);
   U19803 : BUF_X1 port map( A => n25590, Z => n30832);
   U19804 : BUF_X1 port map( A => n25590, Z => n30833);
   U19805 : BUF_X1 port map( A => n25590, Z => n30834);
   U19806 : BUF_X1 port map( A => n25457, Z => n30856);
   U19807 : BUF_X1 port map( A => n25457, Z => n30857);
   U19808 : BUF_X1 port map( A => n25457, Z => n30858);
   U19809 : BUF_X1 port map( A => n25457, Z => n30859);
   U19810 : BUF_X1 port map( A => n25457, Z => n30860);
   U19811 : BUF_X1 port map( A => n25305, Z => n30906);
   U19812 : BUF_X1 port map( A => n25305, Z => n30907);
   U19813 : BUF_X1 port map( A => n25305, Z => n30908);
   U19814 : BUF_X1 port map( A => n25305, Z => n30909);
   U19815 : BUF_X1 port map( A => n25305, Z => n30910);
   U19816 : BUF_X1 port map( A => n25155, Z => n31136);
   U19817 : BUF_X1 port map( A => n30749, Z => n30751);
   U19818 : BUF_X1 port map( A => n30453, Z => n30455);
   U19819 : BUF_X1 port map( A => n30454, Z => n30458);
   U19820 : BUF_X1 port map( A => n30453, Z => n30457);
   U19821 : BUF_X1 port map( A => n30453, Z => n30456);
   U19822 : BUF_X1 port map( A => n30749, Z => n30752);
   U19823 : BUF_X1 port map( A => n30749, Z => n30753);
   U19824 : BUF_X1 port map( A => n30750, Z => n30754);
   U19825 : BUF_X1 port map( A => n30750, Z => n30755);
   U19826 : BUF_X1 port map( A => n25803, Z => n30768);
   U19827 : BUF_X1 port map( A => n25803, Z => n30769);
   U19828 : BUF_X1 port map( A => n25803, Z => n30770);
   U19829 : BUF_X1 port map( A => n25803, Z => n30771);
   U19830 : BUF_X1 port map( A => n25803, Z => n30772);
   U19831 : BUF_X1 port map( A => n26095, Z => n30645);
   U19832 : BUF_X1 port map( A => n26095, Z => n30646);
   U19833 : BUF_X1 port map( A => n26098, Z => n30633);
   U19834 : BUF_X1 port map( A => n26098, Z => n30634);
   U19835 : BUF_X1 port map( A => n26095, Z => n30647);
   U19836 : BUF_X1 port map( A => n26095, Z => n30648);
   U19837 : BUF_X1 port map( A => n26098, Z => n30635);
   U19838 : BUF_X1 port map( A => n26098, Z => n30636);
   U19839 : BUF_X1 port map( A => n26095, Z => n30644);
   U19840 : BUF_X1 port map( A => n26098, Z => n30632);
   U19841 : BUF_X1 port map( A => n26090, Z => n30669);
   U19842 : BUF_X1 port map( A => n26090, Z => n30670);
   U19843 : BUF_X1 port map( A => n26090, Z => n30671);
   U19844 : BUF_X1 port map( A => n26090, Z => n30672);
   U19845 : BUF_X1 port map( A => n26093, Z => n30657);
   U19846 : BUF_X1 port map( A => n26093, Z => n30658);
   U19847 : BUF_X1 port map( A => n26093, Z => n30659);
   U19848 : BUF_X1 port map( A => n26093, Z => n30660);
   U19849 : BUF_X1 port map( A => n26090, Z => n30668);
   U19850 : BUF_X1 port map( A => n26093, Z => n30656);
   U19851 : BUF_X1 port map( A => n25942, Z => n30718);
   U19852 : BUF_X1 port map( A => n26235, Z => n30594);
   U19853 : BUF_X1 port map( A => n26249, Z => n30582);
   U19854 : BUF_X1 port map( A => n26249, Z => n30583);
   U19855 : BUF_X1 port map( A => n26249, Z => n30584);
   U19856 : BUF_X1 port map( A => n26249, Z => n30585);
   U19857 : BUF_X1 port map( A => n26249, Z => n30586);
   U19858 : BUF_X1 port map( A => n26235, Z => n30595);
   U19859 : BUF_X1 port map( A => n26235, Z => n30596);
   U19860 : BUF_X1 port map( A => n26235, Z => n30597);
   U19861 : BUF_X1 port map( A => n26235, Z => n30598);
   U19862 : BUF_X1 port map( A => n25956, Z => n30706);
   U19863 : BUF_X1 port map( A => n25956, Z => n30707);
   U19864 : BUF_X1 port map( A => n25956, Z => n30708);
   U19865 : BUF_X1 port map( A => n25956, Z => n30709);
   U19866 : BUF_X1 port map( A => n25956, Z => n30710);
   U19867 : BUF_X1 port map( A => n25942, Z => n30719);
   U19868 : BUF_X1 port map( A => n25942, Z => n30720);
   U19869 : BUF_X1 port map( A => n25942, Z => n30721);
   U19870 : BUF_X1 port map( A => n25942, Z => n30722);
   U19871 : BUF_X1 port map( A => n25805, Z => n30756);
   U19872 : BUF_X1 port map( A => n25805, Z => n30757);
   U19873 : BUF_X1 port map( A => n25805, Z => n30758);
   U19874 : BUF_X1 port map( A => n25805, Z => n30759);
   U19875 : BUF_X1 port map( A => n25805, Z => n30760);
   U19876 : BUF_X1 port map( A => n25669, Z => n30806);
   U19877 : BUF_X1 port map( A => n25669, Z => n30807);
   U19878 : BUF_X1 port map( A => n25669, Z => n30808);
   U19879 : BUF_X1 port map( A => n25669, Z => n30809);
   U19880 : BUF_X1 port map( A => n25669, Z => n30810);
   U19881 : BUF_X1 port map( A => n25656, Z => n30818);
   U19882 : BUF_X1 port map( A => n25656, Z => n30819);
   U19883 : BUF_X1 port map( A => n25656, Z => n30820);
   U19884 : BUF_X1 port map( A => n25656, Z => n30821);
   U19885 : BUF_X1 port map( A => n25656, Z => n30822);
   U19886 : BUF_X1 port map( A => n25384, Z => n30882);
   U19887 : BUF_X1 port map( A => n25384, Z => n30883);
   U19888 : BUF_X1 port map( A => n25384, Z => n30884);
   U19889 : BUF_X1 port map( A => n25384, Z => n30885);
   U19890 : BUF_X1 port map( A => n25384, Z => n30886);
   U19891 : BUF_X1 port map( A => n25370, Z => n30894);
   U19892 : BUF_X1 port map( A => n25370, Z => n30895);
   U19893 : BUF_X1 port map( A => n25370, Z => n30896);
   U19894 : BUF_X1 port map( A => n25370, Z => n30897);
   U19895 : BUF_X1 port map( A => n25370, Z => n30898);
   U19896 : BUF_X1 port map( A => n25234, Z => n30932);
   U19897 : BUF_X1 port map( A => n25234, Z => n30933);
   U19898 : BUF_X1 port map( A => n25234, Z => n30934);
   U19899 : BUF_X1 port map( A => n25234, Z => n30935);
   U19900 : BUF_X1 port map( A => n25234, Z => n30936);
   U19901 : NAND2_X1 port map( A1 => n31176, A2 => n30851, ZN => n25523);
   U19902 : NAND2_X1 port map( A1 => n31175, A2 => n30801, ZN => n25672);
   U19903 : NAND2_X1 port map( A1 => n31176, A2 => n30927, ZN => n25238);
   U19904 : NAND2_X1 port map( A1 => n31176, A2 => n30877, ZN => n25387);
   U19905 : NAND2_X1 port map( A1 => n31177, A2 => n30564, ZN => n26318);
   U19906 : NAND2_X1 port map( A1 => n31175, A2 => n30751, ZN => n25809);
   U19907 : NAND2_X1 port map( A1 => n31175, A2 => n30701, ZN => n25959);
   U19908 : NAND2_X1 port map( A1 => n31175, A2 => n30688, ZN => n26025);
   U19909 : NAND2_X1 port map( A1 => n31174, A2 => n30627, ZN => n26104);
   U19910 : NAND2_X1 port map( A1 => n31175, A2 => n30577, ZN => n26252);
   U19911 : NAND2_X1 port map( A1 => n31175, A2 => n30614, ZN => n26170);
   U19912 : NAND2_X1 port map( A1 => n31174, A2 => n30738, ZN => n25876);
   U19913 : NAND2_X1 port map( A1 => n31176, A2 => n30788, ZN => n25738);
   U19914 : NAND2_X1 port map( A1 => n31175, A2 => n30838, ZN => n25590);
   U19915 : NAND2_X1 port map( A1 => n31176, A2 => n30864, ZN => n25457);
   U19916 : NAND2_X1 port map( A1 => n31176, A2 => n30914, ZN => n25305);
   U19917 : BUF_X1 port map( A => n30454, Z => n30459);
   U19918 : NAND2_X1 port map( A1 => n31177, A2 => n31142, ZN => n25155);
   U19919 : BUF_X1 port map( A => n25154, Z => n31146);
   U19920 : BUF_X1 port map( A => n30849, Z => n30851);
   U19921 : BUF_X1 port map( A => n30799, Z => n30801);
   U19922 : BUF_X1 port map( A => n30925, Z => n30927);
   U19923 : BUF_X1 port map( A => n30875, Z => n30877);
   U19924 : BUF_X1 port map( A => n30699, Z => n30701);
   U19925 : BUF_X1 port map( A => n30686, Z => n30688);
   U19926 : BUF_X1 port map( A => n30625, Z => n30627);
   U19927 : BUF_X1 port map( A => n30575, Z => n30577);
   U19928 : BUF_X1 port map( A => n30562, Z => n30564);
   U19929 : BUF_X1 port map( A => n30612, Z => n30614);
   U19930 : BUF_X1 port map( A => n30736, Z => n30738);
   U19931 : BUF_X1 port map( A => n30786, Z => n30788);
   U19932 : BUF_X1 port map( A => n30836, Z => n30838);
   U19933 : BUF_X1 port map( A => n30862, Z => n30864);
   U19934 : BUF_X1 port map( A => n30912, Z => n30914);
   U19935 : BUF_X1 port map( A => n30849, Z => n30852);
   U19936 : BUF_X1 port map( A => n30849, Z => n30853);
   U19937 : BUF_X1 port map( A => n30850, Z => n30854);
   U19938 : BUF_X1 port map( A => n30799, Z => n30802);
   U19939 : BUF_X1 port map( A => n30799, Z => n30803);
   U19940 : BUF_X1 port map( A => n30800, Z => n30804);
   U19941 : BUF_X1 port map( A => n30925, Z => n30928);
   U19942 : BUF_X1 port map( A => n30925, Z => n30929);
   U19943 : BUF_X1 port map( A => n30926, Z => n30930);
   U19944 : BUF_X1 port map( A => n30875, Z => n30878);
   U19945 : BUF_X1 port map( A => n30875, Z => n30879);
   U19946 : BUF_X1 port map( A => n30876, Z => n30880);
   U19947 : BUF_X1 port map( A => n30850, Z => n30855);
   U19948 : BUF_X1 port map( A => n30800, Z => n30805);
   U19949 : BUF_X1 port map( A => n30926, Z => n30931);
   U19950 : BUF_X1 port map( A => n30876, Z => n30881);
   U19951 : BUF_X1 port map( A => n30699, Z => n30702);
   U19952 : BUF_X1 port map( A => n30699, Z => n30703);
   U19953 : BUF_X1 port map( A => n30686, Z => n30689);
   U19954 : BUF_X1 port map( A => n30686, Z => n30690);
   U19955 : BUF_X1 port map( A => n30625, Z => n30628);
   U19956 : BUF_X1 port map( A => n30625, Z => n30629);
   U19957 : BUF_X1 port map( A => n30700, Z => n30704);
   U19958 : BUF_X1 port map( A => n30687, Z => n30691);
   U19959 : BUF_X1 port map( A => n30626, Z => n30630);
   U19960 : BUF_X1 port map( A => n30575, Z => n30578);
   U19961 : BUF_X1 port map( A => n30575, Z => n30579);
   U19962 : BUF_X1 port map( A => n30576, Z => n30580);
   U19963 : BUF_X1 port map( A => n30562, Z => n30565);
   U19964 : BUF_X1 port map( A => n30562, Z => n30566);
   U19965 : BUF_X1 port map( A => n30563, Z => n30567);
   U19966 : BUF_X1 port map( A => n30563, Z => n30568);
   U19967 : BUF_X1 port map( A => n30700, Z => n30705);
   U19968 : BUF_X1 port map( A => n30687, Z => n30692);
   U19969 : BUF_X1 port map( A => n30626, Z => n30631);
   U19970 : BUF_X1 port map( A => n30576, Z => n30581);
   U19971 : BUF_X1 port map( A => n30612, Z => n30615);
   U19972 : BUF_X1 port map( A => n30612, Z => n30616);
   U19973 : BUF_X1 port map( A => n30613, Z => n30617);
   U19974 : BUF_X1 port map( A => n30613, Z => n30618);
   U19975 : BUF_X1 port map( A => n30736, Z => n30739);
   U19976 : BUF_X1 port map( A => n30736, Z => n30740);
   U19977 : BUF_X1 port map( A => n30737, Z => n30741);
   U19978 : BUF_X1 port map( A => n30737, Z => n30742);
   U19979 : BUF_X1 port map( A => n30786, Z => n30789);
   U19980 : BUF_X1 port map( A => n30786, Z => n30790);
   U19981 : BUF_X1 port map( A => n30787, Z => n30791);
   U19982 : BUF_X1 port map( A => n30787, Z => n30792);
   U19983 : BUF_X1 port map( A => n30836, Z => n30839);
   U19984 : BUF_X1 port map( A => n30836, Z => n30840);
   U19985 : BUF_X1 port map( A => n30837, Z => n30841);
   U19986 : BUF_X1 port map( A => n30837, Z => n30842);
   U19987 : BUF_X1 port map( A => n30862, Z => n30865);
   U19988 : BUF_X1 port map( A => n30862, Z => n30866);
   U19989 : BUF_X1 port map( A => n30863, Z => n30867);
   U19990 : BUF_X1 port map( A => n30863, Z => n30868);
   U19991 : BUF_X1 port map( A => n30912, Z => n30915);
   U19992 : BUF_X1 port map( A => n30912, Z => n30916);
   U19993 : BUF_X1 port map( A => n30913, Z => n30917);
   U19994 : BUF_X1 port map( A => n30913, Z => n30918);
   U19995 : BUF_X1 port map( A => n25154, Z => n31142);
   U19996 : BUF_X1 port map( A => n25154, Z => n31145);
   U19997 : BUF_X1 port map( A => n25154, Z => n31143);
   U19998 : BUF_X1 port map( A => n25154, Z => n31144);
   U19999 : BUF_X1 port map( A => n28076, Z => n30225);
   U20000 : BUF_X1 port map( A => n28076, Z => n30226);
   U20001 : BUF_X1 port map( A => n28076, Z => n30227);
   U20002 : BUF_X1 port map( A => n28076, Z => n30228);
   U20003 : BUF_X1 port map( A => n28076, Z => n30229);
   U20004 : BUF_X1 port map( A => n31156, Z => n31177);
   U20005 : BUF_X1 port map( A => n31156, Z => n31178);
   U20006 : BUF_X1 port map( A => n31157, Z => n31179);
   U20007 : BUF_X1 port map( A => n31157, Z => n31184);
   U20008 : BUF_X1 port map( A => n31157, Z => n31183);
   U20009 : BUF_X1 port map( A => n31157, Z => n31182);
   U20010 : BUF_X1 port map( A => n31157, Z => n31181);
   U20011 : BUF_X1 port map( A => n31157, Z => n31180);
   U20012 : BUF_X1 port map( A => n31158, Z => n31186);
   U20013 : BUF_X1 port map( A => n31158, Z => n31185);
   U20014 : NAND2_X1 port map( A1 => n31175, A2 => n30774, ZN => n25803);
   U20015 : NAND2_X1 port map( A1 => n31174, A2 => n30674, ZN => n26090);
   U20016 : NAND2_X1 port map( A1 => n31174, A2 => n30638, ZN => n26098);
   U20017 : NAND2_X1 port map( A1 => n31174, A2 => n30662, ZN => n26093);
   U20018 : NAND2_X1 port map( A1 => n31176, A2 => n30650, ZN => n26095);
   U20019 : NAND2_X1 port map( A1 => n31175, A2 => n30588, ZN => n26249);
   U20020 : NAND2_X1 port map( A1 => n31175, A2 => n30600, ZN => n26235);
   U20021 : NAND2_X1 port map( A1 => n31176, A2 => n30712, ZN => n25956);
   U20022 : NAND2_X1 port map( A1 => n31175, A2 => n30724, ZN => n25942);
   U20023 : NAND2_X1 port map( A1 => n31175, A2 => n30762, ZN => n25805);
   U20024 : NAND2_X1 port map( A1 => n31176, A2 => n30812, ZN => n25669);
   U20025 : NAND2_X1 port map( A1 => n31174, A2 => n30824, ZN => n25656);
   U20026 : NAND2_X1 port map( A1 => n31176, A2 => n30888, ZN => n25384);
   U20027 : NAND2_X1 port map( A1 => n31176, A2 => n30900, ZN => n25370);
   U20028 : NAND2_X1 port map( A1 => n31176, A2 => n30938, ZN => n25234);
   U20029 : BUF_X1 port map( A => n31154, Z => n31161);
   U20030 : BUF_X1 port map( A => n31154, Z => n31162);
   U20031 : BUF_X1 port map( A => n31154, Z => n31163);
   U20032 : BUF_X1 port map( A => n31155, Z => n31172);
   U20033 : BUF_X1 port map( A => n31156, Z => n31173);
   U20034 : BUF_X1 port map( A => n31155, Z => n31171);
   U20035 : BUF_X1 port map( A => n31154, Z => n31164);
   U20036 : BUF_X1 port map( A => n31154, Z => n31166);
   U20037 : BUF_X1 port map( A => n31155, Z => n31167);
   U20038 : BUF_X1 port map( A => n31154, Z => n31165);
   U20039 : BUF_X1 port map( A => n31155, Z => n31168);
   U20040 : BUF_X1 port map( A => n31155, Z => n31169);
   U20041 : BUF_X1 port map( A => n31155, Z => n31170);
   U20042 : BUF_X1 port map( A => n31156, Z => n31174);
   U20043 : BUF_X1 port map( A => n31156, Z => n31175);
   U20044 : BUF_X1 port map( A => n31156, Z => n31176);
   U20045 : BUF_X1 port map( A => n25807, Z => n30749);
   U20046 : BUF_X1 port map( A => n26346, Z => n30453);
   U20047 : BUF_X1 port map( A => n25807, Z => n30750);
   U20048 : BUF_X1 port map( A => n26346, Z => n30454);
   U20049 : OAI21_X1 port map( B1 => n25231, B2 => n25232, A => n31163, ZN => 
                           n25154);
   U20050 : BUF_X1 port map( A => n28078, Z => n30213);
   U20051 : BUF_X1 port map( A => n28073, Z => n30237);
   U20052 : BUF_X1 port map( A => n28083, Z => n30189);
   U20053 : BUF_X1 port map( A => n28088, Z => n30165);
   U20054 : BUF_X1 port map( A => n28054, Z => n30309);
   U20055 : BUF_X1 port map( A => n28049, Z => n30333);
   U20056 : BUF_X1 port map( A => n28059, Z => n30285);
   U20057 : BUF_X1 port map( A => n28064, Z => n30261);
   U20058 : BUF_X1 port map( A => n28078, Z => n30214);
   U20059 : BUF_X1 port map( A => n28073, Z => n30238);
   U20060 : BUF_X1 port map( A => n28083, Z => n30190);
   U20061 : BUF_X1 port map( A => n28088, Z => n30166);
   U20062 : BUF_X1 port map( A => n28054, Z => n30310);
   U20063 : BUF_X1 port map( A => n28049, Z => n30334);
   U20064 : BUF_X1 port map( A => n28059, Z => n30286);
   U20065 : BUF_X1 port map( A => n28064, Z => n30262);
   U20066 : BUF_X1 port map( A => n28078, Z => n30215);
   U20067 : BUF_X1 port map( A => n28073, Z => n30239);
   U20068 : BUF_X1 port map( A => n28083, Z => n30191);
   U20069 : BUF_X1 port map( A => n28088, Z => n30167);
   U20070 : BUF_X1 port map( A => n28054, Z => n30311);
   U20071 : BUF_X1 port map( A => n28049, Z => n30335);
   U20072 : BUF_X1 port map( A => n28059, Z => n30287);
   U20073 : BUF_X1 port map( A => n28064, Z => n30263);
   U20074 : BUF_X1 port map( A => n28078, Z => n30216);
   U20075 : BUF_X1 port map( A => n28073, Z => n30240);
   U20076 : BUF_X1 port map( A => n28083, Z => n30192);
   U20077 : BUF_X1 port map( A => n28088, Z => n30168);
   U20078 : BUF_X1 port map( A => n28054, Z => n30312);
   U20079 : BUF_X1 port map( A => n28049, Z => n30336);
   U20080 : BUF_X1 port map( A => n28059, Z => n30288);
   U20081 : BUF_X1 port map( A => n28064, Z => n30264);
   U20082 : BUF_X1 port map( A => n28078, Z => n30217);
   U20083 : BUF_X1 port map( A => n28073, Z => n30241);
   U20084 : BUF_X1 port map( A => n28083, Z => n30193);
   U20085 : BUF_X1 port map( A => n28088, Z => n30169);
   U20086 : BUF_X1 port map( A => n28054, Z => n30313);
   U20087 : BUF_X1 port map( A => n28049, Z => n30337);
   U20088 : BUF_X1 port map( A => n28059, Z => n30289);
   U20089 : BUF_X1 port map( A => n28064, Z => n30265);
   U20090 : BUF_X1 port map( A => n26352, Z => n30441);
   U20091 : BUF_X1 port map( A => n26371, Z => n30369);
   U20092 : BUF_X1 port map( A => n26357, Z => n30417);
   U20093 : BUF_X1 port map( A => n26364, Z => n30393);
   U20094 : BUF_X1 port map( A => n26333, Z => n30514);
   U20095 : BUF_X1 port map( A => n26338, Z => n30490);
   U20096 : BUF_X1 port map( A => n26343, Z => n30466);
   U20097 : BUF_X1 port map( A => n26328, Z => n30538);
   U20098 : BUF_X1 port map( A => n26352, Z => n30442);
   U20099 : BUF_X1 port map( A => n26371, Z => n30370);
   U20100 : BUF_X1 port map( A => n26357, Z => n30418);
   U20101 : BUF_X1 port map( A => n26364, Z => n30394);
   U20102 : BUF_X1 port map( A => n26343, Z => n30467);
   U20103 : BUF_X1 port map( A => n26333, Z => n30515);
   U20104 : BUF_X1 port map( A => n26338, Z => n30491);
   U20105 : BUF_X1 port map( A => n26328, Z => n30539);
   U20106 : BUF_X1 port map( A => n26343, Z => n30468);
   U20107 : BUF_X1 port map( A => n26333, Z => n30516);
   U20108 : BUF_X1 port map( A => n26338, Z => n30492);
   U20109 : BUF_X1 port map( A => n26328, Z => n30540);
   U20110 : BUF_X1 port map( A => n26352, Z => n30443);
   U20111 : BUF_X1 port map( A => n26371, Z => n30371);
   U20112 : BUF_X1 port map( A => n26357, Z => n30419);
   U20113 : BUF_X1 port map( A => n26364, Z => n30395);
   U20114 : BUF_X1 port map( A => n26343, Z => n30469);
   U20115 : BUF_X1 port map( A => n26333, Z => n30517);
   U20116 : BUF_X1 port map( A => n26338, Z => n30493);
   U20117 : BUF_X1 port map( A => n26328, Z => n30541);
   U20118 : BUF_X1 port map( A => n26352, Z => n30444);
   U20119 : BUF_X1 port map( A => n26371, Z => n30372);
   U20120 : BUF_X1 port map( A => n26357, Z => n30420);
   U20121 : BUF_X1 port map( A => n26364, Z => n30396);
   U20122 : BUF_X1 port map( A => n26343, Z => n30470);
   U20123 : BUF_X1 port map( A => n26333, Z => n30518);
   U20124 : BUF_X1 port map( A => n26338, Z => n30494);
   U20125 : BUF_X1 port map( A => n26328, Z => n30542);
   U20126 : BUF_X1 port map( A => n26352, Z => n30445);
   U20127 : BUF_X1 port map( A => n26371, Z => n30373);
   U20128 : BUF_X1 port map( A => n26357, Z => n30421);
   U20129 : BUF_X1 port map( A => n26364, Z => n30397);
   U20130 : BUF_X1 port map( A => n28093, Z => n30144);
   U20131 : BUF_X1 port map( A => n28093, Z => n30145);
   U20132 : BUF_X1 port map( A => n25151, Z => n31151);
   U20133 : BUF_X1 port map( A => n25151, Z => n31152);
   U20134 : BUF_X1 port map( A => n28044, Z => n30339);
   U20135 : BUF_X1 port map( A => n28044, Z => n30340);
   U20136 : BUF_X1 port map( A => n28044, Z => n30341);
   U20137 : BUF_X1 port map( A => n28044, Z => n30342);
   U20138 : BUF_X1 port map( A => n28044, Z => n30343);
   U20139 : BUF_X1 port map( A => n26323, Z => n30544);
   U20140 : BUF_X1 port map( A => n26323, Z => n30545);
   U20141 : BUF_X1 port map( A => n26323, Z => n30546);
   U20142 : BUF_X1 port map( A => n26323, Z => n30547);
   U20143 : BUF_X1 port map( A => n26323, Z => n30548);
   U20144 : BUF_X1 port map( A => n28079, Z => n30207);
   U20145 : BUF_X1 port map( A => n28074, Z => n30231);
   U20146 : BUF_X1 port map( A => n28084, Z => n30183);
   U20147 : BUF_X1 port map( A => n28089, Z => n30159);
   U20148 : BUF_X1 port map( A => n28055, Z => n30303);
   U20149 : BUF_X1 port map( A => n28050, Z => n30327);
   U20150 : BUF_X1 port map( A => n28060, Z => n30279);
   U20151 : BUF_X1 port map( A => n28065, Z => n30255);
   U20152 : BUF_X1 port map( A => n28079, Z => n30208);
   U20153 : BUF_X1 port map( A => n28074, Z => n30232);
   U20154 : BUF_X1 port map( A => n28084, Z => n30184);
   U20155 : BUF_X1 port map( A => n28089, Z => n30160);
   U20156 : BUF_X1 port map( A => n28055, Z => n30304);
   U20157 : BUF_X1 port map( A => n28050, Z => n30328);
   U20158 : BUF_X1 port map( A => n28060, Z => n30280);
   U20159 : BUF_X1 port map( A => n28065, Z => n30256);
   U20160 : BUF_X1 port map( A => n28079, Z => n30209);
   U20161 : BUF_X1 port map( A => n28074, Z => n30233);
   U20162 : BUF_X1 port map( A => n28084, Z => n30185);
   U20163 : BUF_X1 port map( A => n28089, Z => n30161);
   U20164 : BUF_X1 port map( A => n28055, Z => n30305);
   U20165 : BUF_X1 port map( A => n28050, Z => n30329);
   U20166 : BUF_X1 port map( A => n28060, Z => n30281);
   U20167 : BUF_X1 port map( A => n28065, Z => n30257);
   U20168 : BUF_X1 port map( A => n28079, Z => n30210);
   U20169 : BUF_X1 port map( A => n28074, Z => n30234);
   U20170 : BUF_X1 port map( A => n28084, Z => n30186);
   U20171 : BUF_X1 port map( A => n28089, Z => n30162);
   U20172 : BUF_X1 port map( A => n28055, Z => n30306);
   U20173 : BUF_X1 port map( A => n28050, Z => n30330);
   U20174 : BUF_X1 port map( A => n28060, Z => n30282);
   U20175 : BUF_X1 port map( A => n28065, Z => n30258);
   U20176 : BUF_X1 port map( A => n28079, Z => n30211);
   U20177 : BUF_X1 port map( A => n28074, Z => n30235);
   U20178 : BUF_X1 port map( A => n28084, Z => n30187);
   U20179 : BUF_X1 port map( A => n28089, Z => n30163);
   U20180 : BUF_X1 port map( A => n28055, Z => n30307);
   U20181 : BUF_X1 port map( A => n28050, Z => n30331);
   U20182 : BUF_X1 port map( A => n28060, Z => n30283);
   U20183 : BUF_X1 port map( A => n28065, Z => n30259);
   U20184 : BUF_X1 port map( A => n26353, Z => n30435);
   U20185 : BUF_X1 port map( A => n26373, Z => n30363);
   U20186 : BUF_X1 port map( A => n26359, Z => n30411);
   U20187 : BUF_X1 port map( A => n26366, Z => n30387);
   U20188 : BUF_X1 port map( A => n26334, Z => n30508);
   U20189 : BUF_X1 port map( A => n26339, Z => n30484);
   U20190 : BUF_X1 port map( A => n26344, Z => n30460);
   U20191 : BUF_X1 port map( A => n26329, Z => n30532);
   U20192 : BUF_X1 port map( A => n26353, Z => n30436);
   U20193 : BUF_X1 port map( A => n26373, Z => n30364);
   U20194 : BUF_X1 port map( A => n26359, Z => n30412);
   U20195 : BUF_X1 port map( A => n26366, Z => n30388);
   U20196 : BUF_X1 port map( A => n26344, Z => n30461);
   U20197 : BUF_X1 port map( A => n26334, Z => n30509);
   U20198 : BUF_X1 port map( A => n26339, Z => n30485);
   U20199 : BUF_X1 port map( A => n26329, Z => n30533);
   U20200 : BUF_X1 port map( A => n26344, Z => n30462);
   U20201 : BUF_X1 port map( A => n26334, Z => n30510);
   U20202 : BUF_X1 port map( A => n26339, Z => n30486);
   U20203 : BUF_X1 port map( A => n26329, Z => n30534);
   U20204 : BUF_X1 port map( A => n26353, Z => n30437);
   U20205 : BUF_X1 port map( A => n26373, Z => n30365);
   U20206 : BUF_X1 port map( A => n26359, Z => n30413);
   U20207 : BUF_X1 port map( A => n26366, Z => n30389);
   U20208 : BUF_X1 port map( A => n26344, Z => n30463);
   U20209 : BUF_X1 port map( A => n26334, Z => n30511);
   U20210 : BUF_X1 port map( A => n26339, Z => n30487);
   U20211 : BUF_X1 port map( A => n26329, Z => n30535);
   U20212 : BUF_X1 port map( A => n26353, Z => n30438);
   U20213 : BUF_X1 port map( A => n26373, Z => n30366);
   U20214 : BUF_X1 port map( A => n26359, Z => n30414);
   U20215 : BUF_X1 port map( A => n26366, Z => n30390);
   U20216 : BUF_X1 port map( A => n26344, Z => n30464);
   U20217 : BUF_X1 port map( A => n26334, Z => n30512);
   U20218 : BUF_X1 port map( A => n26339, Z => n30488);
   U20219 : BUF_X1 port map( A => n26329, Z => n30536);
   U20220 : BUF_X1 port map( A => n26353, Z => n30439);
   U20221 : BUF_X1 port map( A => n26373, Z => n30367);
   U20222 : BUF_X1 port map( A => n26359, Z => n30415);
   U20223 : BUF_X1 port map( A => n26366, Z => n30391);
   U20224 : BUF_X1 port map( A => n25655, Z => n30828);
   U20225 : BUF_X1 port map( A => n25369, Z => n30904);
   U20226 : BUF_X1 port map( A => n26234, Z => n30604);
   U20227 : BUF_X1 port map( A => n25941, Z => n30728);
   U20228 : BUF_X1 port map( A => n25802, Z => n30774);
   U20229 : BUF_X1 port map( A => n26094, Z => n30650);
   U20230 : BUF_X1 port map( A => n26097, Z => n30638);
   U20231 : BUF_X1 port map( A => n26089, Z => n30674);
   U20232 : BUF_X1 port map( A => n26092, Z => n30662);
   U20233 : BUF_X1 port map( A => n26248, Z => n30588);
   U20234 : BUF_X1 port map( A => n26234, Z => n30600);
   U20235 : BUF_X1 port map( A => n25955, Z => n30712);
   U20236 : BUF_X1 port map( A => n25941, Z => n30724);
   U20237 : BUF_X1 port map( A => n25804, Z => n30762);
   U20238 : BUF_X1 port map( A => n25668, Z => n30812);
   U20239 : BUF_X1 port map( A => n25655, Z => n30824);
   U20240 : BUF_X1 port map( A => n25383, Z => n30888);
   U20241 : BUF_X1 port map( A => n25369, Z => n30900);
   U20242 : BUF_X1 port map( A => n25233, Z => n30938);
   U20243 : BUF_X1 port map( A => n25802, Z => n30775);
   U20244 : BUF_X1 port map( A => n25802, Z => n30776);
   U20245 : BUF_X1 port map( A => n25802, Z => n30777);
   U20246 : BUF_X1 port map( A => n25802, Z => n30778);
   U20247 : BUF_X1 port map( A => n26094, Z => n30652);
   U20248 : BUF_X1 port map( A => n26097, Z => n30640);
   U20249 : BUF_X1 port map( A => n26094, Z => n30653);
   U20250 : BUF_X1 port map( A => n26094, Z => n30654);
   U20251 : BUF_X1 port map( A => n26097, Z => n30641);
   U20252 : BUF_X1 port map( A => n26097, Z => n30642);
   U20253 : BUF_X1 port map( A => n26094, Z => n30651);
   U20254 : BUF_X1 port map( A => n26097, Z => n30639);
   U20255 : BUF_X1 port map( A => n26089, Z => n30676);
   U20256 : BUF_X1 port map( A => n26089, Z => n30677);
   U20257 : BUF_X1 port map( A => n26089, Z => n30678);
   U20258 : BUF_X1 port map( A => n26092, Z => n30664);
   U20259 : BUF_X1 port map( A => n26092, Z => n30665);
   U20260 : BUF_X1 port map( A => n26092, Z => n30666);
   U20261 : BUF_X1 port map( A => n26089, Z => n30675);
   U20262 : BUF_X1 port map( A => n26092, Z => n30663);
   U20263 : BUF_X1 port map( A => n26248, Z => n30589);
   U20264 : BUF_X1 port map( A => n26248, Z => n30590);
   U20265 : BUF_X1 port map( A => n26248, Z => n30591);
   U20266 : BUF_X1 port map( A => n26248, Z => n30592);
   U20267 : BUF_X1 port map( A => n26234, Z => n30603);
   U20268 : BUF_X1 port map( A => n26234, Z => n30601);
   U20269 : BUF_X1 port map( A => n26234, Z => n30602);
   U20270 : BUF_X1 port map( A => n25955, Z => n30713);
   U20271 : BUF_X1 port map( A => n25955, Z => n30714);
   U20272 : BUF_X1 port map( A => n25955, Z => n30715);
   U20273 : BUF_X1 port map( A => n25955, Z => n30716);
   U20274 : BUF_X1 port map( A => n25941, Z => n30727);
   U20275 : BUF_X1 port map( A => n25941, Z => n30725);
   U20276 : BUF_X1 port map( A => n25941, Z => n30726);
   U20277 : BUF_X1 port map( A => n25804, Z => n30763);
   U20278 : BUF_X1 port map( A => n25804, Z => n30764);
   U20279 : BUF_X1 port map( A => n25804, Z => n30765);
   U20280 : BUF_X1 port map( A => n25804, Z => n30766);
   U20281 : BUF_X1 port map( A => n25668, Z => n30813);
   U20282 : BUF_X1 port map( A => n25668, Z => n30814);
   U20283 : BUF_X1 port map( A => n25668, Z => n30815);
   U20284 : BUF_X1 port map( A => n25668, Z => n30816);
   U20285 : BUF_X1 port map( A => n25655, Z => n30827);
   U20286 : BUF_X1 port map( A => n25655, Z => n30825);
   U20287 : BUF_X1 port map( A => n25655, Z => n30826);
   U20288 : BUF_X1 port map( A => n25383, Z => n30889);
   U20289 : BUF_X1 port map( A => n25383, Z => n30890);
   U20290 : BUF_X1 port map( A => n25383, Z => n30891);
   U20291 : BUF_X1 port map( A => n25383, Z => n30892);
   U20292 : BUF_X1 port map( A => n25369, Z => n30903);
   U20293 : BUF_X1 port map( A => n25369, Z => n30901);
   U20294 : BUF_X1 port map( A => n25369, Z => n30902);
   U20295 : BUF_X1 port map( A => n25233, Z => n30939);
   U20296 : BUF_X1 port map( A => n25233, Z => n30940);
   U20297 : BUF_X1 port map( A => n25233, Z => n30941);
   U20298 : BUF_X1 port map( A => n25233, Z => n30942);
   U20299 : BUF_X1 port map( A => n26355, Z => n30429);
   U20300 : BUF_X1 port map( A => n26369, Z => n30381);
   U20301 : BUF_X1 port map( A => n26336, Z => n30502);
   U20302 : BUF_X1 port map( A => n26341, Z => n30478);
   U20303 : BUF_X1 port map( A => n26355, Z => n30430);
   U20304 : BUF_X1 port map( A => n26369, Z => n30382);
   U20305 : BUF_X1 port map( A => n26336, Z => n30503);
   U20306 : BUF_X1 port map( A => n26341, Z => n30479);
   U20307 : BUF_X1 port map( A => n26336, Z => n30504);
   U20308 : BUF_X1 port map( A => n26341, Z => n30480);
   U20309 : BUF_X1 port map( A => n26355, Z => n30431);
   U20310 : BUF_X1 port map( A => n26369, Z => n30383);
   U20311 : BUF_X1 port map( A => n26336, Z => n30505);
   U20312 : BUF_X1 port map( A => n26341, Z => n30481);
   U20313 : BUF_X1 port map( A => n26355, Z => n30432);
   U20314 : BUF_X1 port map( A => n26369, Z => n30384);
   U20315 : BUF_X1 port map( A => n26336, Z => n30506);
   U20316 : BUF_X1 port map( A => n26341, Z => n30482);
   U20317 : BUF_X1 port map( A => n26355, Z => n30433);
   U20318 : BUF_X1 port map( A => n26369, Z => n30385);
   U20319 : BUF_X1 port map( A => n28081, Z => n30201);
   U20320 : BUF_X1 port map( A => n28086, Z => n30177);
   U20321 : BUF_X1 port map( A => n28091, Z => n30153);
   U20322 : BUF_X1 port map( A => n28057, Z => n30297);
   U20323 : BUF_X1 port map( A => n28052, Z => n30321);
   U20324 : BUF_X1 port map( A => n28062, Z => n30273);
   U20325 : BUF_X1 port map( A => n28067, Z => n30249);
   U20326 : BUF_X1 port map( A => n28081, Z => n30202);
   U20327 : BUF_X1 port map( A => n28086, Z => n30178);
   U20328 : BUF_X1 port map( A => n28091, Z => n30154);
   U20329 : BUF_X1 port map( A => n28057, Z => n30298);
   U20330 : BUF_X1 port map( A => n28052, Z => n30322);
   U20331 : BUF_X1 port map( A => n28062, Z => n30274);
   U20332 : BUF_X1 port map( A => n28067, Z => n30250);
   U20333 : BUF_X1 port map( A => n28081, Z => n30203);
   U20334 : BUF_X1 port map( A => n28086, Z => n30179);
   U20335 : BUF_X1 port map( A => n28091, Z => n30155);
   U20336 : BUF_X1 port map( A => n28057, Z => n30299);
   U20337 : BUF_X1 port map( A => n28052, Z => n30323);
   U20338 : BUF_X1 port map( A => n28062, Z => n30275);
   U20339 : BUF_X1 port map( A => n28067, Z => n30251);
   U20340 : BUF_X1 port map( A => n28081, Z => n30204);
   U20341 : BUF_X1 port map( A => n28086, Z => n30180);
   U20342 : BUF_X1 port map( A => n28091, Z => n30156);
   U20343 : BUF_X1 port map( A => n28057, Z => n30300);
   U20344 : BUF_X1 port map( A => n28052, Z => n30324);
   U20345 : BUF_X1 port map( A => n28062, Z => n30276);
   U20346 : BUF_X1 port map( A => n28067, Z => n30252);
   U20347 : BUF_X1 port map( A => n28081, Z => n30205);
   U20348 : BUF_X1 port map( A => n28086, Z => n30181);
   U20349 : BUF_X1 port map( A => n28091, Z => n30157);
   U20350 : BUF_X1 port map( A => n28057, Z => n30301);
   U20351 : BUF_X1 port map( A => n28052, Z => n30325);
   U20352 : BUF_X1 port map( A => n28062, Z => n30277);
   U20353 : BUF_X1 port map( A => n28067, Z => n30253);
   U20354 : BUF_X1 port map( A => n26376, Z => n30357);
   U20355 : BUF_X1 port map( A => n26362, Z => n30405);
   U20356 : BUF_X1 port map( A => n26331, Z => n30526);
   U20357 : BUF_X1 port map( A => n26376, Z => n30358);
   U20358 : BUF_X1 port map( A => n26362, Z => n30406);
   U20359 : BUF_X1 port map( A => n26331, Z => n30527);
   U20360 : BUF_X1 port map( A => n26331, Z => n30528);
   U20361 : BUF_X1 port map( A => n26376, Z => n30359);
   U20362 : BUF_X1 port map( A => n26362, Z => n30407);
   U20363 : BUF_X1 port map( A => n26331, Z => n30529);
   U20364 : BUF_X1 port map( A => n26376, Z => n30360);
   U20365 : BUF_X1 port map( A => n26362, Z => n30408);
   U20366 : BUF_X1 port map( A => n26331, Z => n30530);
   U20367 : BUF_X1 port map( A => n26376, Z => n30361);
   U20368 : BUF_X1 port map( A => n26362, Z => n30409);
   U20369 : NAND2_X1 port map( A1 => n29300, A2 => n29287, ZN => n28076);
   U20370 : BUF_X1 port map( A => n26370, Z => n30375);
   U20371 : BUF_X1 port map( A => n26337, Z => n30496);
   U20372 : BUF_X1 port map( A => n26342, Z => n30472);
   U20373 : BUF_X1 port map( A => n26370, Z => n30376);
   U20374 : BUF_X1 port map( A => n26337, Z => n30497);
   U20375 : BUF_X1 port map( A => n26342, Z => n30473);
   U20376 : BUF_X1 port map( A => n26337, Z => n30498);
   U20377 : BUF_X1 port map( A => n26342, Z => n30474);
   U20378 : BUF_X1 port map( A => n26370, Z => n30377);
   U20379 : BUF_X1 port map( A => n26337, Z => n30499);
   U20380 : BUF_X1 port map( A => n26342, Z => n30475);
   U20381 : BUF_X1 port map( A => n26370, Z => n30378);
   U20382 : BUF_X1 port map( A => n26337, Z => n30500);
   U20383 : BUF_X1 port map( A => n26342, Z => n30476);
   U20384 : BUF_X1 port map( A => n26370, Z => n30379);
   U20385 : BUF_X1 port map( A => n28082, Z => n30195);
   U20386 : BUF_X1 port map( A => n28077, Z => n30219);
   U20387 : BUF_X1 port map( A => n28087, Z => n30171);
   U20388 : BUF_X1 port map( A => n28092, Z => n30147);
   U20389 : BUF_X1 port map( A => n28058, Z => n30291);
   U20390 : BUF_X1 port map( A => n28053, Z => n30315);
   U20391 : BUF_X1 port map( A => n28063, Z => n30267);
   U20392 : BUF_X1 port map( A => n28068, Z => n30243);
   U20393 : BUF_X1 port map( A => n28082, Z => n30196);
   U20394 : BUF_X1 port map( A => n28077, Z => n30220);
   U20395 : BUF_X1 port map( A => n28087, Z => n30172);
   U20396 : BUF_X1 port map( A => n28092, Z => n30148);
   U20397 : BUF_X1 port map( A => n28058, Z => n30292);
   U20398 : BUF_X1 port map( A => n28053, Z => n30316);
   U20399 : BUF_X1 port map( A => n28063, Z => n30268);
   U20400 : BUF_X1 port map( A => n28068, Z => n30244);
   U20401 : BUF_X1 port map( A => n28082, Z => n30197);
   U20402 : BUF_X1 port map( A => n28077, Z => n30221);
   U20403 : BUF_X1 port map( A => n28087, Z => n30173);
   U20404 : BUF_X1 port map( A => n28092, Z => n30149);
   U20405 : BUF_X1 port map( A => n28058, Z => n30293);
   U20406 : BUF_X1 port map( A => n28053, Z => n30317);
   U20407 : BUF_X1 port map( A => n28063, Z => n30269);
   U20408 : BUF_X1 port map( A => n28068, Z => n30245);
   U20409 : BUF_X1 port map( A => n28082, Z => n30198);
   U20410 : BUF_X1 port map( A => n28077, Z => n30222);
   U20411 : BUF_X1 port map( A => n28087, Z => n30174);
   U20412 : BUF_X1 port map( A => n28092, Z => n30150);
   U20413 : BUF_X1 port map( A => n28058, Z => n30294);
   U20414 : BUF_X1 port map( A => n28053, Z => n30318);
   U20415 : BUF_X1 port map( A => n28063, Z => n30270);
   U20416 : BUF_X1 port map( A => n28068, Z => n30246);
   U20417 : BUF_X1 port map( A => n28082, Z => n30199);
   U20418 : BUF_X1 port map( A => n28077, Z => n30223);
   U20419 : BUF_X1 port map( A => n28087, Z => n30175);
   U20420 : BUF_X1 port map( A => n28092, Z => n30151);
   U20421 : BUF_X1 port map( A => n28058, Z => n30295);
   U20422 : BUF_X1 port map( A => n28053, Z => n30319);
   U20423 : BUF_X1 port map( A => n28063, Z => n30271);
   U20424 : BUF_X1 port map( A => n28068, Z => n30247);
   U20425 : BUF_X1 port map( A => n26356, Z => n30423);
   U20426 : BUF_X1 port map( A => n26377, Z => n30351);
   U20427 : BUF_X1 port map( A => n26363, Z => n30399);
   U20428 : BUF_X1 port map( A => n26347, Z => n30447);
   U20429 : BUF_X1 port map( A => n26332, Z => n30520);
   U20430 : BUF_X1 port map( A => n26356, Z => n30424);
   U20431 : BUF_X1 port map( A => n26377, Z => n30352);
   U20432 : BUF_X1 port map( A => n26363, Z => n30400);
   U20433 : BUF_X1 port map( A => n26347, Z => n30448);
   U20434 : BUF_X1 port map( A => n26332, Z => n30521);
   U20435 : BUF_X1 port map( A => n26347, Z => n30449);
   U20436 : BUF_X1 port map( A => n26332, Z => n30522);
   U20437 : BUF_X1 port map( A => n26356, Z => n30425);
   U20438 : BUF_X1 port map( A => n26377, Z => n30353);
   U20439 : BUF_X1 port map( A => n26363, Z => n30401);
   U20440 : BUF_X1 port map( A => n26347, Z => n30450);
   U20441 : BUF_X1 port map( A => n26332, Z => n30523);
   U20442 : BUF_X1 port map( A => n26356, Z => n30426);
   U20443 : BUF_X1 port map( A => n26377, Z => n30354);
   U20444 : BUF_X1 port map( A => n26363, Z => n30402);
   U20445 : BUF_X1 port map( A => n26347, Z => n30451);
   U20446 : BUF_X1 port map( A => n26332, Z => n30524);
   U20447 : BUF_X1 port map( A => n26356, Z => n30427);
   U20448 : BUF_X1 port map( A => n26377, Z => n30355);
   U20449 : BUF_X1 port map( A => n26363, Z => n30403);
   U20450 : BUF_X1 port map( A => n28093, Z => n30141);
   U20451 : BUF_X1 port map( A => n28093, Z => n30142);
   U20452 : BUF_X1 port map( A => n28093, Z => n30143);
   U20453 : BUF_X1 port map( A => n25151, Z => n31148);
   U20454 : BUF_X1 port map( A => n25151, Z => n31149);
   U20455 : BUF_X1 port map( A => n25151, Z => n31150);
   U20456 : OAI21_X1 port map( B1 => n25232, B2 => n25873, A => n31162, ZN => 
                           n25807);
   U20457 : BUF_X1 port map( A => n31159, Z => n31156);
   U20458 : BUF_X1 port map( A => n31159, Z => n31157);
   U20459 : BUF_X1 port map( A => n31160, Z => n31154);
   U20460 : BUF_X1 port map( A => n31160, Z => n31155);
   U20461 : NAND2_X1 port map( A1 => n28013, A2 => n28006, ZN => n26346);
   U20462 : BUF_X1 port map( A => n25455, Z => n30862);
   U20463 : BUF_X1 port map( A => n25303, Z => n30912);
   U20464 : BUF_X1 port map( A => n25236, Z => n30925);
   U20465 : BUF_X1 port map( A => n25385, Z => n30875);
   U20466 : BUF_X1 port map( A => n25521, Z => n30849);
   U20467 : BUF_X1 port map( A => n25670, Z => n30799);
   U20468 : BUF_X1 port map( A => n25736, Z => n30786);
   U20469 : BUF_X1 port map( A => n25588, Z => n30836);
   U20470 : BUF_X1 port map( A => n25957, Z => n30699);
   U20471 : BUF_X1 port map( A => n26023, Z => n30686);
   U20472 : BUF_X1 port map( A => n26102, Z => n30625);
   U20473 : BUF_X1 port map( A => n26250, Z => n30575);
   U20474 : BUF_X1 port map( A => n26316, Z => n30562);
   U20475 : BUF_X1 port map( A => n26168, Z => n30612);
   U20476 : BUF_X1 port map( A => n25874, Z => n30736);
   U20477 : BUF_X1 port map( A => n31159, Z => n31158);
   U20478 : BUF_X1 port map( A => n25455, Z => n30863);
   U20479 : BUF_X1 port map( A => n25303, Z => n30913);
   U20480 : BUF_X1 port map( A => n25236, Z => n30926);
   U20481 : BUF_X1 port map( A => n25385, Z => n30876);
   U20482 : BUF_X1 port map( A => n25521, Z => n30850);
   U20483 : BUF_X1 port map( A => n25670, Z => n30800);
   U20484 : BUF_X1 port map( A => n25736, Z => n30787);
   U20485 : BUF_X1 port map( A => n25588, Z => n30837);
   U20486 : BUF_X1 port map( A => n26316, Z => n30563);
   U20487 : BUF_X1 port map( A => n25957, Z => n30700);
   U20488 : BUF_X1 port map( A => n26023, Z => n30687);
   U20489 : BUF_X1 port map( A => n26102, Z => n30626);
   U20490 : BUF_X1 port map( A => n26250, Z => n30576);
   U20491 : BUF_X1 port map( A => n26168, Z => n30613);
   U20492 : BUF_X1 port map( A => n25874, Z => n30737);
   U20493 : NOR2_X1 port map( A1 => n29305, A2 => n29308, ZN => n29287);
   U20494 : OAI21_X1 port map( B1 => n25235, B2 => n25382, A => n31162, ZN => 
                           n25383);
   U20495 : OAI21_X1 port map( B1 => n25451, B2 => n25587, A => n31162, ZN => 
                           n25802);
   U20496 : OAI21_X1 port map( B1 => n25302, B2 => n25587, A => n31163, ZN => 
                           n25655);
   U20497 : OAI21_X1 port map( B1 => n25451, B2 => n25654, A => n31162, ZN => 
                           n25804);
   U20498 : OAI21_X1 port map( B1 => n25302, B2 => n25654, A => n31163, ZN => 
                           n25668);
   U20499 : OAI21_X1 port map( B1 => n25451, B2 => n25873, A => n31162, ZN => 
                           n26089);
   U20500 : OAI21_X1 port map( B1 => n25232, B2 => n26099, A => n31161, ZN => 
                           n26097);
   U20501 : OAI21_X1 port map( B1 => n25451, B2 => n25940, A => n31162, ZN => 
                           n26092);
   U20502 : OAI21_X1 port map( B1 => n25232, B2 => n26096, A => n31162, ZN => 
                           n26094);
   U20503 : OAI21_X1 port map( B1 => n25382, B2 => n26099, A => n31161, ZN => 
                           n26248);
   U20504 : OAI21_X1 port map( B1 => n25382, B2 => n26096, A => n31161, ZN => 
                           n26234);
   U20505 : OAI21_X1 port map( B1 => n25302, B2 => n25940, A => n31161, ZN => 
                           n25955);
   U20506 : OAI21_X1 port map( B1 => n25302, B2 => n25873, A => n31162, ZN => 
                           n25941);
   U20507 : OAI21_X1 port map( B1 => n25231, B2 => n25382, A => n31163, ZN => 
                           n25369);
   U20508 : OAI21_X1 port map( B1 => n25232, B2 => n25235, A => n31162, ZN => 
                           n25233);
   U20509 : NOR3_X1 port map( A1 => n29288, A2 => n29306, A3 => n29293, ZN => 
                           n29300);
   U20510 : NOR2_X1 port map( A1 => n28028, A2 => n28033, ZN => n28006);
   U20511 : NOR3_X1 port map( A1 => n28024, A2 => n28029, A3 => n28007, ZN => 
                           n28013);
   U20512 : BUF_X1 port map( A => n28040, Z => n30345);
   U20513 : BUF_X1 port map( A => n28040, Z => n30346);
   U20514 : BUF_X1 port map( A => n28040, Z => n30347);
   U20515 : BUF_X1 port map( A => n28040, Z => n30348);
   U20516 : BUF_X1 port map( A => n28040, Z => n30349);
   U20517 : BUF_X1 port map( A => n26319, Z => n30550);
   U20518 : BUF_X1 port map( A => n26319, Z => n30551);
   U20519 : BUF_X1 port map( A => n26319, Z => n30552);
   U20520 : BUF_X1 port map( A => n26319, Z => n30553);
   U20521 : BUF_X1 port map( A => n26319, Z => n30554);
   U20522 : OAI21_X1 port map( B1 => n25152, B2 => n29313, A => n31161, ZN => 
                           n28093);
   U20523 : OAI21_X1 port map( B1 => n25152, B2 => n25153, A => n31162, ZN => 
                           n25151);
   U20524 : NAND2_X1 port map( A1 => n26100, A2 => n26101, ZN => n25232);
   U20525 : NAND2_X1 port map( A1 => n28005, A2 => n28019, ZN => n26356);
   U20526 : NAND2_X1 port map( A1 => n29286, A2 => n29302, ZN => n28082);
   U20527 : NAND2_X1 port map( A1 => n29286, A2 => n29300, ZN => n28086);
   U20528 : NAND2_X1 port map( A1 => n29286, A2 => n29299, ZN => n28087);
   U20529 : NAND2_X1 port map( A1 => n29287, A2 => n29299, ZN => n28077);
   U20530 : BUF_X1 port map( A => n25230, Z => n30944);
   U20531 : BUF_X1 port map( A => n25228, Z => n30947);
   U20532 : BUF_X1 port map( A => n25226, Z => n30950);
   U20533 : BUF_X1 port map( A => n25224, Z => n30953);
   U20534 : BUF_X1 port map( A => n25222, Z => n30956);
   U20535 : BUF_X1 port map( A => n25220, Z => n30959);
   U20536 : BUF_X1 port map( A => n25218, Z => n30962);
   U20537 : BUF_X1 port map( A => n25216, Z => n30965);
   U20538 : BUF_X1 port map( A => n25214, Z => n30968);
   U20539 : BUF_X1 port map( A => n25212, Z => n30971);
   U20540 : BUF_X1 port map( A => n25210, Z => n30974);
   U20541 : BUF_X1 port map( A => n25208, Z => n30977);
   U20542 : BUF_X1 port map( A => n25207, Z => n30980);
   U20543 : BUF_X1 port map( A => n25206, Z => n30983);
   U20544 : BUF_X1 port map( A => n25205, Z => n30986);
   U20545 : BUF_X1 port map( A => n25204, Z => n30989);
   U20546 : BUF_X1 port map( A => n25203, Z => n30992);
   U20547 : BUF_X1 port map( A => n25202, Z => n30995);
   U20548 : BUF_X1 port map( A => n25201, Z => n30998);
   U20549 : BUF_X1 port map( A => n25200, Z => n31001);
   U20550 : BUF_X1 port map( A => n25199, Z => n31004);
   U20551 : BUF_X1 port map( A => n25198, Z => n31007);
   U20552 : BUF_X1 port map( A => n25197, Z => n31010);
   U20553 : BUF_X1 port map( A => n25196, Z => n31013);
   U20554 : BUF_X1 port map( A => n25195, Z => n31016);
   U20555 : BUF_X1 port map( A => n25194, Z => n31019);
   U20556 : BUF_X1 port map( A => n25193, Z => n31022);
   U20557 : BUF_X1 port map( A => n25192, Z => n31025);
   U20558 : BUF_X1 port map( A => n25191, Z => n31028);
   U20559 : BUF_X1 port map( A => n25190, Z => n31031);
   U20560 : BUF_X1 port map( A => n25189, Z => n31034);
   U20561 : BUF_X1 port map( A => n25188, Z => n31037);
   U20562 : BUF_X1 port map( A => n25187, Z => n31040);
   U20563 : BUF_X1 port map( A => n25186, Z => n31043);
   U20564 : BUF_X1 port map( A => n25185, Z => n31046);
   U20565 : BUF_X1 port map( A => n25184, Z => n31049);
   U20566 : BUF_X1 port map( A => n25183, Z => n31052);
   U20567 : BUF_X1 port map( A => n25182, Z => n31055);
   U20568 : BUF_X1 port map( A => n25181, Z => n31058);
   U20569 : BUF_X1 port map( A => n25180, Z => n31061);
   U20570 : BUF_X1 port map( A => n25179, Z => n31064);
   U20571 : BUF_X1 port map( A => n25178, Z => n31067);
   U20572 : BUF_X1 port map( A => n25177, Z => n31070);
   U20573 : BUF_X1 port map( A => n25176, Z => n31073);
   U20574 : BUF_X1 port map( A => n25175, Z => n31076);
   U20575 : BUF_X1 port map( A => n25174, Z => n31079);
   U20576 : BUF_X1 port map( A => n25173, Z => n31082);
   U20577 : BUF_X1 port map( A => n25172, Z => n31085);
   U20578 : BUF_X1 port map( A => n25171, Z => n31088);
   U20579 : BUF_X1 port map( A => n25170, Z => n31091);
   U20580 : BUF_X1 port map( A => n25169, Z => n31094);
   U20581 : BUF_X1 port map( A => n25168, Z => n31097);
   U20582 : BUF_X1 port map( A => n25167, Z => n31100);
   U20583 : BUF_X1 port map( A => n25166, Z => n31103);
   U20584 : BUF_X1 port map( A => n25165, Z => n31106);
   U20585 : BUF_X1 port map( A => n25164, Z => n31109);
   U20586 : BUF_X1 port map( A => n25163, Z => n31112);
   U20587 : BUF_X1 port map( A => n25162, Z => n31115);
   U20588 : BUF_X1 port map( A => n25161, Z => n31118);
   U20589 : BUF_X1 port map( A => n25160, Z => n31121);
   U20590 : BUF_X1 port map( A => n25159, Z => n31124);
   U20591 : BUF_X1 port map( A => n25158, Z => n31127);
   U20592 : BUF_X1 port map( A => n25157, Z => n31130);
   U20593 : BUF_X1 port map( A => n25156, Z => n31133);
   U20594 : NAND2_X1 port map( A1 => n28003, A2 => n28019, ZN => n26377);
   U20595 : NAND2_X1 port map( A1 => n28003, A2 => n28020, ZN => n26376);
   U20596 : NAND2_X1 port map( A1 => n28003, A2 => n28009, ZN => n26363);
   U20597 : BUF_X1 port map( A => n25230, Z => n30945);
   U20598 : BUF_X1 port map( A => n25228, Z => n30948);
   U20599 : BUF_X1 port map( A => n25226, Z => n30951);
   U20600 : BUF_X1 port map( A => n25224, Z => n30954);
   U20601 : BUF_X1 port map( A => n25222, Z => n30957);
   U20602 : BUF_X1 port map( A => n25220, Z => n30960);
   U20603 : BUF_X1 port map( A => n25218, Z => n30963);
   U20604 : BUF_X1 port map( A => n25216, Z => n30966);
   U20605 : BUF_X1 port map( A => n25214, Z => n30969);
   U20606 : BUF_X1 port map( A => n25212, Z => n30972);
   U20607 : BUF_X1 port map( A => n25210, Z => n30975);
   U20608 : BUF_X1 port map( A => n25208, Z => n30978);
   U20609 : BUF_X1 port map( A => n25207, Z => n30981);
   U20610 : BUF_X1 port map( A => n25206, Z => n30984);
   U20611 : BUF_X1 port map( A => n25205, Z => n30987);
   U20612 : BUF_X1 port map( A => n25204, Z => n30990);
   U20613 : BUF_X1 port map( A => n25203, Z => n30993);
   U20614 : BUF_X1 port map( A => n25202, Z => n30996);
   U20615 : BUF_X1 port map( A => n25201, Z => n30999);
   U20616 : BUF_X1 port map( A => n25200, Z => n31002);
   U20617 : BUF_X1 port map( A => n25199, Z => n31005);
   U20618 : BUF_X1 port map( A => n25198, Z => n31008);
   U20619 : BUF_X1 port map( A => n25197, Z => n31011);
   U20620 : BUF_X1 port map( A => n25196, Z => n31014);
   U20621 : BUF_X1 port map( A => n25195, Z => n31017);
   U20622 : BUF_X1 port map( A => n25194, Z => n31020);
   U20623 : BUF_X1 port map( A => n25193, Z => n31023);
   U20624 : BUF_X1 port map( A => n25192, Z => n31026);
   U20625 : BUF_X1 port map( A => n25191, Z => n31029);
   U20626 : BUF_X1 port map( A => n25190, Z => n31032);
   U20627 : BUF_X1 port map( A => n25189, Z => n31035);
   U20628 : BUF_X1 port map( A => n25188, Z => n31038);
   U20629 : BUF_X1 port map( A => n25187, Z => n31041);
   U20630 : BUF_X1 port map( A => n25186, Z => n31044);
   U20631 : BUF_X1 port map( A => n25185, Z => n31047);
   U20632 : BUF_X1 port map( A => n25184, Z => n31050);
   U20633 : BUF_X1 port map( A => n25183, Z => n31053);
   U20634 : BUF_X1 port map( A => n25182, Z => n31056);
   U20635 : BUF_X1 port map( A => n25181, Z => n31059);
   U20636 : BUF_X1 port map( A => n25180, Z => n31062);
   U20637 : BUF_X1 port map( A => n25179, Z => n31065);
   U20638 : BUF_X1 port map( A => n25178, Z => n31068);
   U20639 : BUF_X1 port map( A => n25177, Z => n31071);
   U20640 : BUF_X1 port map( A => n25176, Z => n31074);
   U20641 : BUF_X1 port map( A => n25175, Z => n31077);
   U20642 : BUF_X1 port map( A => n25174, Z => n31080);
   U20643 : BUF_X1 port map( A => n25173, Z => n31083);
   U20644 : BUF_X1 port map( A => n25172, Z => n31086);
   U20645 : BUF_X1 port map( A => n25171, Z => n31089);
   U20646 : BUF_X1 port map( A => n25170, Z => n31092);
   U20647 : BUF_X1 port map( A => n25169, Z => n31095);
   U20648 : BUF_X1 port map( A => n25168, Z => n31098);
   U20649 : BUF_X1 port map( A => n25167, Z => n31101);
   U20650 : BUF_X1 port map( A => n25166, Z => n31104);
   U20651 : BUF_X1 port map( A => n25165, Z => n31107);
   U20652 : BUF_X1 port map( A => n25164, Z => n31110);
   U20653 : BUF_X1 port map( A => n25163, Z => n31113);
   U20654 : BUF_X1 port map( A => n25162, Z => n31116);
   U20655 : BUF_X1 port map( A => n25161, Z => n31119);
   U20656 : BUF_X1 port map( A => n25160, Z => n31122);
   U20657 : BUF_X1 port map( A => n25159, Z => n31125);
   U20658 : BUF_X1 port map( A => n25158, Z => n31128);
   U20659 : BUF_X1 port map( A => n25157, Z => n31131);
   U20660 : BUF_X1 port map( A => n25156, Z => n31134);
   U20661 : NAND2_X1 port map( A1 => n28020, A2 => n28005, ZN => n26355);
   U20662 : NAND2_X1 port map( A1 => n29302, A2 => n29284, ZN => n28092);
   U20663 : NAND2_X1 port map( A1 => n28009, A2 => n28005, ZN => n26342);
   U20664 : NAND2_X1 port map( A1 => n28002, A2 => n28005, ZN => n26336);
   U20665 : NAND2_X1 port map( A1 => n28000, A2 => n28005, ZN => n26337);
   U20666 : NAND2_X1 port map( A1 => n28010, A2 => n28005, ZN => n26341);
   U20667 : NAND2_X1 port map( A1 => n28013, A2 => n28005, ZN => n26369);
   U20668 : NAND2_X1 port map( A1 => n28012, A2 => n28005, ZN => n26370);
   U20669 : NAND2_X1 port map( A1 => n29303, A2 => n29286, ZN => n28081);
   U20670 : NAND2_X1 port map( A1 => n29303, A2 => n29284, ZN => n28091);
   U20671 : NAND2_X1 port map( A1 => n28010, A2 => n28003, ZN => n26362);
   U20672 : NAND2_X1 port map( A1 => n29283, A2 => n29282, ZN => n28052);
   U20673 : NAND2_X1 port map( A1 => n29281, A2 => n29282, ZN => n28053);
   U20674 : NAND2_X1 port map( A1 => n28002, A2 => n28001, ZN => n26331);
   U20675 : NAND2_X1 port map( A1 => n28000, A2 => n28001, ZN => n26332);
   U20676 : NAND2_X1 port map( A1 => n29283, A2 => n29286, ZN => n28057);
   U20677 : NAND2_X1 port map( A1 => n29281, A2 => n29286, ZN => n28058);
   U20678 : NAND2_X1 port map( A1 => n29291, A2 => n29287, ZN => n28062);
   U20679 : NAND2_X1 port map( A1 => n29290, A2 => n29287, ZN => n28063);
   U20680 : NAND2_X1 port map( A1 => n29291, A2 => n29284, ZN => n28067);
   U20681 : NAND2_X1 port map( A1 => n29290, A2 => n29284, ZN => n28068);
   U20682 : NAND2_X1 port map( A1 => n28012, A2 => n28006, ZN => n26347);
   U20683 : OAI22_X1 port map( A1 => n30805, A2 => n25675, B1 => n31125, B2 => 
                           n30798, ZN => n7109);
   U20684 : OAI22_X1 port map( A1 => n30805, A2 => n25674, B1 => n31128, B2 => 
                           n30798, ZN => n7110);
   U20685 : OAI22_X1 port map( A1 => n30805, A2 => n25673, B1 => n31131, B2 => 
                           n30798, ZN => n7111);
   U20686 : OAI22_X1 port map( A1 => n30805, A2 => n25671, B1 => n31134, B2 => 
                           n30798, ZN => n7112);
   U20687 : OAI22_X1 port map( A1 => n30568, A2 => n26430, B1 => n31124, B2 => 
                           n30561, ZN => n5890);
   U20688 : OAI22_X1 port map( A1 => n30568, A2 => n26404, B1 => n31127, B2 => 
                           n30561, ZN => n5892);
   U20689 : OAI22_X1 port map( A1 => n30568, A2 => n26378, B1 => n31130, B2 => 
                           n30561, ZN => n5894);
   U20690 : OAI22_X1 port map( A1 => n30568, A2 => n26317, B1 => n31133, B2 => 
                           n30561, ZN => n5896);
   U20691 : OAI22_X1 port map( A1 => n30705, A2 => n25962, B1 => n31125, B2 => 
                           n30698, ZN => n6597);
   U20692 : OAI22_X1 port map( A1 => n30705, A2 => n25961, B1 => n31128, B2 => 
                           n30698, ZN => n6598);
   U20693 : OAI22_X1 port map( A1 => n30705, A2 => n25960, B1 => n31131, B2 => 
                           n30698, ZN => n6599);
   U20694 : OAI22_X1 port map( A1 => n30705, A2 => n25958, B1 => n31134, B2 => 
                           n30698, ZN => n6600);
   U20695 : OAI22_X1 port map( A1 => n30692, A2 => n26028, B1 => n31125, B2 => 
                           n30685, ZN => n6533);
   U20696 : OAI22_X1 port map( A1 => n30692, A2 => n26027, B1 => n31128, B2 => 
                           n30685, ZN => n6534);
   U20697 : OAI22_X1 port map( A1 => n30692, A2 => n26026, B1 => n31131, B2 => 
                           n30685, ZN => n6535);
   U20698 : OAI22_X1 port map( A1 => n30692, A2 => n26024, B1 => n31134, B2 => 
                           n30685, ZN => n6536);
   U20699 : OAI22_X1 port map( A1 => n30581, A2 => n26255, B1 => n31126, B2 => 
                           n30574, ZN => n5957);
   U20700 : OAI22_X1 port map( A1 => n30581, A2 => n26254, B1 => n31129, B2 => 
                           n30574, ZN => n5958);
   U20701 : OAI22_X1 port map( A1 => n30581, A2 => n26253, B1 => n31132, B2 => 
                           n30574, ZN => n5959);
   U20702 : OAI22_X1 port map( A1 => n30581, A2 => n26251, B1 => n31135, B2 => 
                           n30574, ZN => n5960);
   U20703 : OAI22_X1 port map( A1 => n30792, A2 => n25741, B1 => n31125, B2 => 
                           n30785, ZN => n7045);
   U20704 : OAI22_X1 port map( A1 => n30792, A2 => n25740, B1 => n31128, B2 => 
                           n30785, ZN => n7046);
   U20705 : OAI22_X1 port map( A1 => n30792, A2 => n25739, B1 => n31131, B2 => 
                           n30785, ZN => n7047);
   U20706 : OAI22_X1 port map( A1 => n30792, A2 => n25737, B1 => n31134, B2 => 
                           n30785, ZN => n7048);
   U20707 : OAI22_X1 port map( A1 => n30578, A2 => n26303, B1 => n30982, B2 => 
                           n30570, ZN => n5909);
   U20708 : OAI22_X1 port map( A1 => n30578, A2 => n26302, B1 => n30985, B2 => 
                           n30570, ZN => n5910);
   U20709 : OAI22_X1 port map( A1 => n30578, A2 => n26301, B1 => n30988, B2 => 
                           n30570, ZN => n5911);
   U20710 : OAI22_X1 port map( A1 => n30578, A2 => n26300, B1 => n30991, B2 => 
                           n30570, ZN => n5912);
   U20711 : OAI22_X1 port map( A1 => n30578, A2 => n26299, B1 => n30994, B2 => 
                           n30570, ZN => n5913);
   U20712 : OAI22_X1 port map( A1 => n30578, A2 => n26298, B1 => n30997, B2 => 
                           n30570, ZN => n5914);
   U20713 : OAI22_X1 port map( A1 => n30578, A2 => n26297, B1 => n31000, B2 => 
                           n30570, ZN => n5915);
   U20714 : OAI22_X1 port map( A1 => n30578, A2 => n26296, B1 => n31003, B2 => 
                           n30570, ZN => n5916);
   U20715 : OAI22_X1 port map( A1 => n30578, A2 => n26295, B1 => n31006, B2 => 
                           n30570, ZN => n5917);
   U20716 : OAI22_X1 port map( A1 => n30578, A2 => n26294, B1 => n31009, B2 => 
                           n30570, ZN => n5918);
   U20717 : OAI22_X1 port map( A1 => n30578, A2 => n26293, B1 => n31012, B2 => 
                           n30570, ZN => n5919);
   U20718 : OAI22_X1 port map( A1 => n30578, A2 => n26292, B1 => n31015, B2 => 
                           n30570, ZN => n5920);
   U20719 : OAI22_X1 port map( A1 => n30578, A2 => n26291, B1 => n31018, B2 => 
                           n30571, ZN => n5921);
   U20720 : OAI22_X1 port map( A1 => n30579, A2 => n26290, B1 => n31021, B2 => 
                           n30571, ZN => n5922);
   U20721 : OAI22_X1 port map( A1 => n30579, A2 => n26289, B1 => n31024, B2 => 
                           n30571, ZN => n5923);
   U20722 : OAI22_X1 port map( A1 => n30579, A2 => n26288, B1 => n31027, B2 => 
                           n30571, ZN => n5924);
   U20723 : OAI22_X1 port map( A1 => n30579, A2 => n26287, B1 => n31030, B2 => 
                           n30571, ZN => n5925);
   U20724 : OAI22_X1 port map( A1 => n30579, A2 => n26286, B1 => n31033, B2 => 
                           n30571, ZN => n5926);
   U20725 : OAI22_X1 port map( A1 => n30579, A2 => n26285, B1 => n31036, B2 => 
                           n30571, ZN => n5927);
   U20726 : OAI22_X1 port map( A1 => n30579, A2 => n26284, B1 => n31039, B2 => 
                           n30571, ZN => n5928);
   U20727 : OAI22_X1 port map( A1 => n30579, A2 => n26283, B1 => n31042, B2 => 
                           n30571, ZN => n5929);
   U20728 : OAI22_X1 port map( A1 => n30579, A2 => n26282, B1 => n31045, B2 => 
                           n30571, ZN => n5930);
   U20729 : OAI22_X1 port map( A1 => n30579, A2 => n26281, B1 => n31048, B2 => 
                           n30571, ZN => n5931);
   U20730 : OAI22_X1 port map( A1 => n30579, A2 => n26280, B1 => n31051, B2 => 
                           n30571, ZN => n5932);
   U20731 : OAI22_X1 port map( A1 => n30579, A2 => n26279, B1 => n31054, B2 => 
                           n30572, ZN => n5933);
   U20732 : OAI22_X1 port map( A1 => n30579, A2 => n26278, B1 => n31057, B2 => 
                           n30572, ZN => n5934);
   U20733 : OAI22_X1 port map( A1 => n30580, A2 => n26277, B1 => n31060, B2 => 
                           n30572, ZN => n5935);
   U20734 : OAI22_X1 port map( A1 => n30580, A2 => n26276, B1 => n31063, B2 => 
                           n30572, ZN => n5936);
   U20735 : OAI22_X1 port map( A1 => n30580, A2 => n26275, B1 => n31066, B2 => 
                           n30572, ZN => n5937);
   U20736 : OAI22_X1 port map( A1 => n30580, A2 => n26274, B1 => n31069, B2 => 
                           n30572, ZN => n5938);
   U20737 : OAI22_X1 port map( A1 => n30580, A2 => n26273, B1 => n31072, B2 => 
                           n30572, ZN => n5939);
   U20738 : OAI22_X1 port map( A1 => n30580, A2 => n26272, B1 => n31075, B2 => 
                           n30572, ZN => n5940);
   U20739 : OAI22_X1 port map( A1 => n30580, A2 => n26271, B1 => n31078, B2 => 
                           n30572, ZN => n5941);
   U20740 : OAI22_X1 port map( A1 => n30580, A2 => n26270, B1 => n31081, B2 => 
                           n30572, ZN => n5942);
   U20741 : OAI22_X1 port map( A1 => n30580, A2 => n26269, B1 => n31084, B2 => 
                           n30572, ZN => n5943);
   U20742 : OAI22_X1 port map( A1 => n30580, A2 => n26268, B1 => n31087, B2 => 
                           n30572, ZN => n5944);
   U20743 : OAI22_X1 port map( A1 => n30580, A2 => n26267, B1 => n31090, B2 => 
                           n30573, ZN => n5945);
   U20744 : OAI22_X1 port map( A1 => n30580, A2 => n26266, B1 => n31093, B2 => 
                           n30573, ZN => n5946);
   U20745 : OAI22_X1 port map( A1 => n30580, A2 => n26265, B1 => n31096, B2 => 
                           n30573, ZN => n5947);
   U20746 : OAI22_X1 port map( A1 => n30581, A2 => n26264, B1 => n31099, B2 => 
                           n30573, ZN => n5948);
   U20747 : OAI22_X1 port map( A1 => n30581, A2 => n26263, B1 => n31102, B2 => 
                           n30573, ZN => n5949);
   U20748 : OAI22_X1 port map( A1 => n30581, A2 => n26262, B1 => n31105, B2 => 
                           n30573, ZN => n5950);
   U20749 : OAI22_X1 port map( A1 => n30581, A2 => n26261, B1 => n31108, B2 => 
                           n30573, ZN => n5951);
   U20750 : OAI22_X1 port map( A1 => n30581, A2 => n26260, B1 => n31111, B2 => 
                           n30573, ZN => n5952);
   U20751 : OAI22_X1 port map( A1 => n30581, A2 => n26259, B1 => n31114, B2 => 
                           n30573, ZN => n5953);
   U20752 : OAI22_X1 port map( A1 => n30581, A2 => n26258, B1 => n31117, B2 => 
                           n30573, ZN => n5954);
   U20753 : OAI22_X1 port map( A1 => n30581, A2 => n26257, B1 => n31120, B2 => 
                           n30573, ZN => n5955);
   U20754 : OAI22_X1 port map( A1 => n30581, A2 => n26256, B1 => n31123, B2 => 
                           n30573, ZN => n5956);
   U20755 : OAI22_X1 port map( A1 => n30577, A2 => n26315, B1 => n30946, B2 => 
                           n30569, ZN => n5897);
   U20756 : OAI22_X1 port map( A1 => n30577, A2 => n26314, B1 => n30949, B2 => 
                           n30569, ZN => n5898);
   U20757 : OAI22_X1 port map( A1 => n30577, A2 => n26313, B1 => n30952, B2 => 
                           n30569, ZN => n5899);
   U20758 : OAI22_X1 port map( A1 => n30577, A2 => n26312, B1 => n30955, B2 => 
                           n30569, ZN => n5900);
   U20759 : OAI22_X1 port map( A1 => n30577, A2 => n26311, B1 => n30958, B2 => 
                           n30569, ZN => n5901);
   U20760 : OAI22_X1 port map( A1 => n30577, A2 => n26310, B1 => n30961, B2 => 
                           n30569, ZN => n5902);
   U20761 : OAI22_X1 port map( A1 => n30577, A2 => n26309, B1 => n30964, B2 => 
                           n30569, ZN => n5903);
   U20762 : OAI22_X1 port map( A1 => n30577, A2 => n26308, B1 => n30967, B2 => 
                           n30569, ZN => n5904);
   U20763 : OAI22_X1 port map( A1 => n30577, A2 => n26307, B1 => n30970, B2 => 
                           n30569, ZN => n5905);
   U20764 : OAI22_X1 port map( A1 => n30577, A2 => n26306, B1 => n30973, B2 => 
                           n30569, ZN => n5906);
   U20765 : OAI22_X1 port map( A1 => n30577, A2 => n26305, B1 => n30976, B2 => 
                           n30569, ZN => n5907);
   U20766 : OAI22_X1 port map( A1 => n30577, A2 => n26304, B1 => n30979, B2 => 
                           n30569, ZN => n5908);
   U20767 : OAI22_X1 port map( A1 => n30604, A2 => n26243, B1 => n30958, B2 => 
                           n30594, ZN => n6029);
   U20768 : OAI22_X1 port map( A1 => n30604, A2 => n26242, B1 => n30961, B2 => 
                           n30594, ZN => n6030);
   U20769 : OAI22_X1 port map( A1 => n30604, A2 => n26241, B1 => n30964, B2 => 
                           n30594, ZN => n6031);
   U20770 : OAI22_X1 port map( A1 => n30604, A2 => n26240, B1 => n30967, B2 => 
                           n30594, ZN => n6032);
   U20771 : OAI22_X1 port map( A1 => n30604, A2 => n26239, B1 => n30970, B2 => 
                           n30594, ZN => n6033);
   U20772 : OAI22_X1 port map( A1 => n30604, A2 => n26238, B1 => n30973, B2 => 
                           n30594, ZN => n6034);
   U20773 : OAI22_X1 port map( A1 => n30604, A2 => n26237, B1 => n30976, B2 => 
                           n30594, ZN => n6035);
   U20774 : OAI22_X1 port map( A1 => n30604, A2 => n26236, B1 => n30979, B2 => 
                           n30594, ZN => n6036);
   U20775 : OAI22_X1 port map( A1 => n30605, A2 => n26247, B1 => n30946, B2 => 
                           n30594, ZN => n6025);
   U20776 : OAI22_X1 port map( A1 => n30605, A2 => n26246, B1 => n30949, B2 => 
                           n30594, ZN => n6026);
   U20777 : OAI22_X1 port map( A1 => n30605, A2 => n26245, B1 => n30952, B2 => 
                           n30594, ZN => n6027);
   U20778 : OAI22_X1 port map( A1 => n30605, A2 => n26244, B1 => n30955, B2 => 
                           n30594, ZN => n6028);
   U20779 : BUF_X1 port map( A => n25230, Z => n30946);
   U20780 : BUF_X1 port map( A => n25228, Z => n30949);
   U20781 : BUF_X1 port map( A => n25226, Z => n30952);
   U20782 : BUF_X1 port map( A => n25224, Z => n30955);
   U20783 : BUF_X1 port map( A => n25222, Z => n30958);
   U20784 : BUF_X1 port map( A => n25220, Z => n30961);
   U20785 : BUF_X1 port map( A => n25218, Z => n30964);
   U20786 : BUF_X1 port map( A => n25216, Z => n30967);
   U20787 : BUF_X1 port map( A => n25214, Z => n30970);
   U20788 : BUF_X1 port map( A => n25212, Z => n30973);
   U20789 : BUF_X1 port map( A => n25210, Z => n30976);
   U20790 : BUF_X1 port map( A => n25208, Z => n30979);
   U20791 : BUF_X1 port map( A => n25207, Z => n30982);
   U20792 : BUF_X1 port map( A => n25206, Z => n30985);
   U20793 : BUF_X1 port map( A => n25205, Z => n30988);
   U20794 : BUF_X1 port map( A => n25204, Z => n30991);
   U20795 : BUF_X1 port map( A => n25203, Z => n30994);
   U20796 : BUF_X1 port map( A => n25202, Z => n30997);
   U20797 : BUF_X1 port map( A => n25201, Z => n31000);
   U20798 : BUF_X1 port map( A => n25200, Z => n31003);
   U20799 : BUF_X1 port map( A => n25199, Z => n31006);
   U20800 : BUF_X1 port map( A => n25198, Z => n31009);
   U20801 : BUF_X1 port map( A => n25197, Z => n31012);
   U20802 : BUF_X1 port map( A => n25196, Z => n31015);
   U20803 : BUF_X1 port map( A => n25195, Z => n31018);
   U20804 : BUF_X1 port map( A => n25194, Z => n31021);
   U20805 : BUF_X1 port map( A => n25193, Z => n31024);
   U20806 : BUF_X1 port map( A => n25192, Z => n31027);
   U20807 : BUF_X1 port map( A => n25191, Z => n31030);
   U20808 : BUF_X1 port map( A => n25190, Z => n31033);
   U20809 : BUF_X1 port map( A => n25189, Z => n31036);
   U20810 : BUF_X1 port map( A => n25188, Z => n31039);
   U20811 : BUF_X1 port map( A => n25187, Z => n31042);
   U20812 : BUF_X1 port map( A => n25186, Z => n31045);
   U20813 : BUF_X1 port map( A => n25185, Z => n31048);
   U20814 : BUF_X1 port map( A => n25184, Z => n31051);
   U20815 : BUF_X1 port map( A => n25183, Z => n31054);
   U20816 : BUF_X1 port map( A => n25182, Z => n31057);
   U20817 : BUF_X1 port map( A => n25181, Z => n31060);
   U20818 : BUF_X1 port map( A => n25180, Z => n31063);
   U20819 : BUF_X1 port map( A => n25179, Z => n31066);
   U20820 : BUF_X1 port map( A => n25178, Z => n31069);
   U20821 : BUF_X1 port map( A => n25177, Z => n31072);
   U20822 : BUF_X1 port map( A => n25176, Z => n31075);
   U20823 : BUF_X1 port map( A => n25175, Z => n31078);
   U20824 : BUF_X1 port map( A => n25174, Z => n31081);
   U20825 : BUF_X1 port map( A => n25173, Z => n31084);
   U20826 : BUF_X1 port map( A => n25172, Z => n31087);
   U20827 : BUF_X1 port map( A => n25171, Z => n31090);
   U20828 : BUF_X1 port map( A => n25170, Z => n31093);
   U20829 : BUF_X1 port map( A => n25169, Z => n31096);
   U20830 : BUF_X1 port map( A => n25168, Z => n31099);
   U20831 : BUF_X1 port map( A => n25167, Z => n31102);
   U20832 : BUF_X1 port map( A => n25166, Z => n31105);
   U20833 : BUF_X1 port map( A => n25165, Z => n31108);
   U20834 : BUF_X1 port map( A => n25164, Z => n31111);
   U20835 : BUF_X1 port map( A => n25163, Z => n31114);
   U20836 : BUF_X1 port map( A => n25162, Z => n31117);
   U20837 : BUF_X1 port map( A => n25161, Z => n31120);
   U20838 : BUF_X1 port map( A => n25160, Z => n31123);
   U20839 : BUF_X1 port map( A => n25159, Z => n31126);
   U20840 : BUF_X1 port map( A => n25158, Z => n31129);
   U20841 : BUF_X1 port map( A => n25157, Z => n31132);
   U20842 : BUF_X1 port map( A => n25156, Z => n31135);
   U20843 : OAI22_X1 port map( A1 => n30801, A2 => n25735, B1 => n30945, B2 => 
                           n30793, ZN => n7049);
   U20844 : OAI22_X1 port map( A1 => n30801, A2 => n25734, B1 => n30948, B2 => 
                           n30793, ZN => n7050);
   U20845 : OAI22_X1 port map( A1 => n30801, A2 => n25733, B1 => n30951, B2 => 
                           n30793, ZN => n7051);
   U20846 : OAI22_X1 port map( A1 => n30801, A2 => n25732, B1 => n30954, B2 => 
                           n30793, ZN => n7052);
   U20847 : OAI22_X1 port map( A1 => n30801, A2 => n25731, B1 => n30957, B2 => 
                           n30793, ZN => n7053);
   U20848 : OAI22_X1 port map( A1 => n30801, A2 => n25730, B1 => n30960, B2 => 
                           n30793, ZN => n7054);
   U20849 : OAI22_X1 port map( A1 => n30801, A2 => n25729, B1 => n30963, B2 => 
                           n30793, ZN => n7055);
   U20850 : OAI22_X1 port map( A1 => n30801, A2 => n25728, B1 => n30966, B2 => 
                           n30793, ZN => n7056);
   U20851 : OAI22_X1 port map( A1 => n30801, A2 => n25727, B1 => n30969, B2 => 
                           n30793, ZN => n7057);
   U20852 : OAI22_X1 port map( A1 => n30801, A2 => n25726, B1 => n30972, B2 => 
                           n30793, ZN => n7058);
   U20853 : OAI22_X1 port map( A1 => n30801, A2 => n25725, B1 => n30975, B2 => 
                           n30793, ZN => n7059);
   U20854 : OAI22_X1 port map( A1 => n30801, A2 => n25724, B1 => n30978, B2 => 
                           n30793, ZN => n7060);
   U20855 : OAI22_X1 port map( A1 => n30802, A2 => n25723, B1 => n30981, B2 => 
                           n30794, ZN => n7061);
   U20856 : OAI22_X1 port map( A1 => n30802, A2 => n25722, B1 => n30984, B2 => 
                           n30794, ZN => n7062);
   U20857 : OAI22_X1 port map( A1 => n30802, A2 => n25721, B1 => n30987, B2 => 
                           n30794, ZN => n7063);
   U20858 : OAI22_X1 port map( A1 => n30802, A2 => n25720, B1 => n30990, B2 => 
                           n30794, ZN => n7064);
   U20859 : OAI22_X1 port map( A1 => n30802, A2 => n25719, B1 => n30993, B2 => 
                           n30794, ZN => n7065);
   U20860 : OAI22_X1 port map( A1 => n30802, A2 => n25718, B1 => n30996, B2 => 
                           n30794, ZN => n7066);
   U20861 : OAI22_X1 port map( A1 => n30802, A2 => n25717, B1 => n30999, B2 => 
                           n30794, ZN => n7067);
   U20862 : OAI22_X1 port map( A1 => n30802, A2 => n25716, B1 => n31002, B2 => 
                           n30794, ZN => n7068);
   U20863 : OAI22_X1 port map( A1 => n30802, A2 => n25715, B1 => n31005, B2 => 
                           n30794, ZN => n7069);
   U20864 : OAI22_X1 port map( A1 => n30802, A2 => n25714, B1 => n31008, B2 => 
                           n30794, ZN => n7070);
   U20865 : OAI22_X1 port map( A1 => n30802, A2 => n25713, B1 => n31011, B2 => 
                           n30794, ZN => n7071);
   U20866 : OAI22_X1 port map( A1 => n30802, A2 => n25712, B1 => n31014, B2 => 
                           n30794, ZN => n7072);
   U20867 : OAI22_X1 port map( A1 => n30802, A2 => n25711, B1 => n31017, B2 => 
                           n30795, ZN => n7073);
   U20868 : OAI22_X1 port map( A1 => n30803, A2 => n25710, B1 => n31020, B2 => 
                           n30795, ZN => n7074);
   U20869 : OAI22_X1 port map( A1 => n30803, A2 => n25709, B1 => n31023, B2 => 
                           n30795, ZN => n7075);
   U20870 : OAI22_X1 port map( A1 => n30803, A2 => n25708, B1 => n31026, B2 => 
                           n30795, ZN => n7076);
   U20871 : OAI22_X1 port map( A1 => n30803, A2 => n25707, B1 => n31029, B2 => 
                           n30795, ZN => n7077);
   U20872 : OAI22_X1 port map( A1 => n30803, A2 => n25706, B1 => n31032, B2 => 
                           n30795, ZN => n7078);
   U20873 : OAI22_X1 port map( A1 => n30803, A2 => n25705, B1 => n31035, B2 => 
                           n30795, ZN => n7079);
   U20874 : OAI22_X1 port map( A1 => n30803, A2 => n25704, B1 => n31038, B2 => 
                           n30795, ZN => n7080);
   U20875 : OAI22_X1 port map( A1 => n30803, A2 => n25703, B1 => n31041, B2 => 
                           n30795, ZN => n7081);
   U20876 : OAI22_X1 port map( A1 => n30803, A2 => n25702, B1 => n31044, B2 => 
                           n30795, ZN => n7082);
   U20877 : OAI22_X1 port map( A1 => n30803, A2 => n25701, B1 => n31047, B2 => 
                           n30795, ZN => n7083);
   U20878 : OAI22_X1 port map( A1 => n30803, A2 => n25700, B1 => n31050, B2 => 
                           n30795, ZN => n7084);
   U20879 : OAI22_X1 port map( A1 => n30803, A2 => n25699, B1 => n31053, B2 => 
                           n30796, ZN => n7085);
   U20880 : OAI22_X1 port map( A1 => n30803, A2 => n25698, B1 => n31056, B2 => 
                           n30796, ZN => n7086);
   U20881 : OAI22_X1 port map( A1 => n30804, A2 => n25697, B1 => n31059, B2 => 
                           n30796, ZN => n7087);
   U20882 : OAI22_X1 port map( A1 => n30804, A2 => n25696, B1 => n31062, B2 => 
                           n30796, ZN => n7088);
   U20883 : OAI22_X1 port map( A1 => n30804, A2 => n25695, B1 => n31065, B2 => 
                           n30796, ZN => n7089);
   U20884 : OAI22_X1 port map( A1 => n30804, A2 => n25694, B1 => n31068, B2 => 
                           n30796, ZN => n7090);
   U20885 : OAI22_X1 port map( A1 => n30804, A2 => n25693, B1 => n31071, B2 => 
                           n30796, ZN => n7091);
   U20886 : OAI22_X1 port map( A1 => n30804, A2 => n25692, B1 => n31074, B2 => 
                           n30796, ZN => n7092);
   U20887 : OAI22_X1 port map( A1 => n30804, A2 => n25691, B1 => n31077, B2 => 
                           n30796, ZN => n7093);
   U20888 : OAI22_X1 port map( A1 => n30804, A2 => n25690, B1 => n31080, B2 => 
                           n30796, ZN => n7094);
   U20889 : OAI22_X1 port map( A1 => n30804, A2 => n25689, B1 => n31083, B2 => 
                           n30796, ZN => n7095);
   U20890 : OAI22_X1 port map( A1 => n30804, A2 => n25688, B1 => n31086, B2 => 
                           n30796, ZN => n7096);
   U20891 : OAI22_X1 port map( A1 => n30804, A2 => n25687, B1 => n31089, B2 => 
                           n30797, ZN => n7097);
   U20892 : OAI22_X1 port map( A1 => n30804, A2 => n25686, B1 => n31092, B2 => 
                           n30797, ZN => n7098);
   U20893 : OAI22_X1 port map( A1 => n30804, A2 => n25685, B1 => n31095, B2 => 
                           n30797, ZN => n7099);
   U20894 : OAI22_X1 port map( A1 => n30805, A2 => n25684, B1 => n31098, B2 => 
                           n30797, ZN => n7100);
   U20895 : OAI22_X1 port map( A1 => n30805, A2 => n25683, B1 => n31101, B2 => 
                           n30797, ZN => n7101);
   U20896 : OAI22_X1 port map( A1 => n30805, A2 => n25682, B1 => n31104, B2 => 
                           n30797, ZN => n7102);
   U20897 : OAI22_X1 port map( A1 => n30805, A2 => n25681, B1 => n31107, B2 => 
                           n30797, ZN => n7103);
   U20898 : OAI22_X1 port map( A1 => n30805, A2 => n25680, B1 => n31110, B2 => 
                           n30797, ZN => n7104);
   U20899 : OAI22_X1 port map( A1 => n30805, A2 => n25679, B1 => n31113, B2 => 
                           n30797, ZN => n7105);
   U20900 : OAI22_X1 port map( A1 => n30805, A2 => n25678, B1 => n31116, B2 => 
                           n30797, ZN => n7106);
   U20901 : OAI22_X1 port map( A1 => n30805, A2 => n25677, B1 => n31119, B2 => 
                           n30797, ZN => n7107);
   U20902 : OAI22_X1 port map( A1 => n30805, A2 => n25676, B1 => n31122, B2 => 
                           n30797, ZN => n7108);
   U20903 : OAI22_X1 port map( A1 => n30829, A2 => n25667, B1 => n30944, B2 => 
                           n30818, ZN => n7177);
   U20904 : OAI22_X1 port map( A1 => n30829, A2 => n25666, B1 => n30947, B2 => 
                           n30818, ZN => n7178);
   U20905 : OAI22_X1 port map( A1 => n30829, A2 => n25665, B1 => n30950, B2 => 
                           n30818, ZN => n7179);
   U20906 : OAI22_X1 port map( A1 => n30829, A2 => n25664, B1 => n30953, B2 => 
                           n30818, ZN => n7180);
   U20907 : OAI22_X1 port map( A1 => n30828, A2 => n25663, B1 => n30956, B2 => 
                           n30818, ZN => n7181);
   U20908 : OAI22_X1 port map( A1 => n30828, A2 => n25662, B1 => n30959, B2 => 
                           n30818, ZN => n7182);
   U20909 : OAI22_X1 port map( A1 => n30828, A2 => n25661, B1 => n30962, B2 => 
                           n30818, ZN => n7183);
   U20910 : OAI22_X1 port map( A1 => n30828, A2 => n25660, B1 => n30965, B2 => 
                           n30818, ZN => n7184);
   U20911 : OAI22_X1 port map( A1 => n30828, A2 => n25659, B1 => n30968, B2 => 
                           n30818, ZN => n7185);
   U20912 : OAI22_X1 port map( A1 => n30828, A2 => n25658, B1 => n30971, B2 => 
                           n30818, ZN => n7186);
   U20913 : OAI22_X1 port map( A1 => n30828, A2 => n25657, B1 => n30974, B2 => 
                           n30818, ZN => n7187);
   U20914 : OAI22_X1 port map( A1 => n30905, A2 => n25381, B1 => n30944, B2 => 
                           n30894, ZN => n7561);
   U20915 : OAI22_X1 port map( A1 => n30905, A2 => n25380, B1 => n30947, B2 => 
                           n30894, ZN => n7562);
   U20916 : OAI22_X1 port map( A1 => n30905, A2 => n25379, B1 => n30950, B2 => 
                           n30894, ZN => n7563);
   U20917 : OAI22_X1 port map( A1 => n30905, A2 => n25378, B1 => n30953, B2 => 
                           n30894, ZN => n7564);
   U20918 : OAI22_X1 port map( A1 => n30904, A2 => n25377, B1 => n30956, B2 => 
                           n30894, ZN => n7565);
   U20919 : OAI22_X1 port map( A1 => n30904, A2 => n25376, B1 => n30959, B2 => 
                           n30894, ZN => n7566);
   U20920 : OAI22_X1 port map( A1 => n30904, A2 => n25375, B1 => n30962, B2 => 
                           n30894, ZN => n7567);
   U20921 : OAI22_X1 port map( A1 => n30904, A2 => n25374, B1 => n30965, B2 => 
                           n30894, ZN => n7568);
   U20922 : OAI22_X1 port map( A1 => n30904, A2 => n25373, B1 => n30968, B2 => 
                           n30894, ZN => n7569);
   U20923 : OAI22_X1 port map( A1 => n30904, A2 => n25372, B1 => n30971, B2 => 
                           n30894, ZN => n7570);
   U20924 : OAI22_X1 port map( A1 => n30904, A2 => n25371, B1 => n30974, B2 => 
                           n30894, ZN => n7571);
   U20925 : OAI22_X1 port map( A1 => n31147, A2 => n25229, B1 => n31136, B2 => 
                           n30944, ZN => n7817);
   U20926 : OAI22_X1 port map( A1 => n31147, A2 => n25227, B1 => n31136, B2 => 
                           n30947, ZN => n7818);
   U20927 : OAI22_X1 port map( A1 => n31147, A2 => n25225, B1 => n31136, B2 => 
                           n30950, ZN => n7819);
   U20928 : OAI22_X1 port map( A1 => n31147, A2 => n25223, B1 => n31136, B2 => 
                           n30953, ZN => n7820);
   U20929 : OAI22_X1 port map( A1 => n31146, A2 => n25221, B1 => n31136, B2 => 
                           n30956, ZN => n7821);
   U20930 : OAI22_X1 port map( A1 => n31146, A2 => n25219, B1 => n31136, B2 => 
                           n30959, ZN => n7822);
   U20931 : OAI22_X1 port map( A1 => n31146, A2 => n25217, B1 => n31136, B2 => 
                           n30962, ZN => n7823);
   U20932 : OAI22_X1 port map( A1 => n31146, A2 => n25215, B1 => n31136, B2 => 
                           n30965, ZN => n7824);
   U20933 : OAI22_X1 port map( A1 => n31146, A2 => n25213, B1 => n31136, B2 => 
                           n30968, ZN => n7825);
   U20934 : OAI22_X1 port map( A1 => n31146, A2 => n25211, B1 => n31136, B2 => 
                           n30971, ZN => n7826);
   U20935 : OAI22_X1 port map( A1 => n31146, A2 => n25209, B1 => n31136, B2 => 
                           n30974, ZN => n7827);
   U20936 : OAI22_X1 port map( A1 => n30702, A2 => n26010, B1 => n30981, B2 => 
                           n30694, ZN => n6549);
   U20937 : OAI22_X1 port map( A1 => n30702, A2 => n26009, B1 => n30984, B2 => 
                           n30694, ZN => n6550);
   U20938 : OAI22_X1 port map( A1 => n30702, A2 => n26008, B1 => n30987, B2 => 
                           n30694, ZN => n6551);
   U20939 : OAI22_X1 port map( A1 => n30702, A2 => n26007, B1 => n30990, B2 => 
                           n30694, ZN => n6552);
   U20940 : OAI22_X1 port map( A1 => n30702, A2 => n26006, B1 => n30993, B2 => 
                           n30694, ZN => n6553);
   U20941 : OAI22_X1 port map( A1 => n30702, A2 => n26005, B1 => n30996, B2 => 
                           n30694, ZN => n6554);
   U20942 : OAI22_X1 port map( A1 => n30702, A2 => n26004, B1 => n30999, B2 => 
                           n30694, ZN => n6555);
   U20943 : OAI22_X1 port map( A1 => n30702, A2 => n26003, B1 => n31002, B2 => 
                           n30694, ZN => n6556);
   U20944 : OAI22_X1 port map( A1 => n30702, A2 => n26002, B1 => n31005, B2 => 
                           n30694, ZN => n6557);
   U20945 : OAI22_X1 port map( A1 => n30702, A2 => n26001, B1 => n31008, B2 => 
                           n30694, ZN => n6558);
   U20946 : OAI22_X1 port map( A1 => n30702, A2 => n26000, B1 => n31011, B2 => 
                           n30694, ZN => n6559);
   U20947 : OAI22_X1 port map( A1 => n30702, A2 => n25999, B1 => n31014, B2 => 
                           n30694, ZN => n6560);
   U20948 : OAI22_X1 port map( A1 => n30702, A2 => n25998, B1 => n31017, B2 => 
                           n30695, ZN => n6561);
   U20949 : OAI22_X1 port map( A1 => n30703, A2 => n25997, B1 => n31020, B2 => 
                           n30695, ZN => n6562);
   U20950 : OAI22_X1 port map( A1 => n30703, A2 => n25996, B1 => n31023, B2 => 
                           n30695, ZN => n6563);
   U20951 : OAI22_X1 port map( A1 => n30703, A2 => n25995, B1 => n31026, B2 => 
                           n30695, ZN => n6564);
   U20952 : OAI22_X1 port map( A1 => n30703, A2 => n25994, B1 => n31029, B2 => 
                           n30695, ZN => n6565);
   U20953 : OAI22_X1 port map( A1 => n30703, A2 => n25993, B1 => n31032, B2 => 
                           n30695, ZN => n6566);
   U20954 : OAI22_X1 port map( A1 => n30703, A2 => n25992, B1 => n31035, B2 => 
                           n30695, ZN => n6567);
   U20955 : OAI22_X1 port map( A1 => n30703, A2 => n25991, B1 => n31038, B2 => 
                           n30695, ZN => n6568);
   U20956 : OAI22_X1 port map( A1 => n30703, A2 => n25990, B1 => n31041, B2 => 
                           n30695, ZN => n6569);
   U20957 : OAI22_X1 port map( A1 => n30703, A2 => n25989, B1 => n31044, B2 => 
                           n30695, ZN => n6570);
   U20958 : OAI22_X1 port map( A1 => n30703, A2 => n25988, B1 => n31047, B2 => 
                           n30695, ZN => n6571);
   U20959 : OAI22_X1 port map( A1 => n30703, A2 => n25987, B1 => n31050, B2 => 
                           n30695, ZN => n6572);
   U20960 : OAI22_X1 port map( A1 => n30703, A2 => n25986, B1 => n31053, B2 => 
                           n30696, ZN => n6573);
   U20961 : OAI22_X1 port map( A1 => n30703, A2 => n25985, B1 => n31056, B2 => 
                           n30696, ZN => n6574);
   U20962 : OAI22_X1 port map( A1 => n30689, A2 => n26076, B1 => n30981, B2 => 
                           n30681, ZN => n6485);
   U20963 : OAI22_X1 port map( A1 => n30689, A2 => n26075, B1 => n30984, B2 => 
                           n30681, ZN => n6486);
   U20964 : OAI22_X1 port map( A1 => n30689, A2 => n26074, B1 => n30987, B2 => 
                           n30681, ZN => n6487);
   U20965 : OAI22_X1 port map( A1 => n30689, A2 => n26073, B1 => n30990, B2 => 
                           n30681, ZN => n6488);
   U20966 : OAI22_X1 port map( A1 => n30689, A2 => n26072, B1 => n30993, B2 => 
                           n30681, ZN => n6489);
   U20967 : OAI22_X1 port map( A1 => n30689, A2 => n26071, B1 => n30996, B2 => 
                           n30681, ZN => n6490);
   U20968 : OAI22_X1 port map( A1 => n30689, A2 => n26070, B1 => n30999, B2 => 
                           n30681, ZN => n6491);
   U20969 : OAI22_X1 port map( A1 => n30689, A2 => n26069, B1 => n31002, B2 => 
                           n30681, ZN => n6492);
   U20970 : OAI22_X1 port map( A1 => n30689, A2 => n26068, B1 => n31005, B2 => 
                           n30681, ZN => n6493);
   U20971 : OAI22_X1 port map( A1 => n30689, A2 => n26067, B1 => n31008, B2 => 
                           n30681, ZN => n6494);
   U20972 : OAI22_X1 port map( A1 => n30689, A2 => n26066, B1 => n31011, B2 => 
                           n30681, ZN => n6495);
   U20973 : OAI22_X1 port map( A1 => n30689, A2 => n26065, B1 => n31014, B2 => 
                           n30681, ZN => n6496);
   U20974 : OAI22_X1 port map( A1 => n30689, A2 => n26064, B1 => n31017, B2 => 
                           n30682, ZN => n6497);
   U20975 : OAI22_X1 port map( A1 => n30690, A2 => n26063, B1 => n31020, B2 => 
                           n30682, ZN => n6498);
   U20976 : OAI22_X1 port map( A1 => n30690, A2 => n26062, B1 => n31023, B2 => 
                           n30682, ZN => n6499);
   U20977 : OAI22_X1 port map( A1 => n30690, A2 => n26061, B1 => n31026, B2 => 
                           n30682, ZN => n6500);
   U20978 : OAI22_X1 port map( A1 => n30690, A2 => n26060, B1 => n31029, B2 => 
                           n30682, ZN => n6501);
   U20979 : OAI22_X1 port map( A1 => n30690, A2 => n26059, B1 => n31032, B2 => 
                           n30682, ZN => n6502);
   U20980 : OAI22_X1 port map( A1 => n30690, A2 => n26058, B1 => n31035, B2 => 
                           n30682, ZN => n6503);
   U20981 : OAI22_X1 port map( A1 => n30690, A2 => n26057, B1 => n31038, B2 => 
                           n30682, ZN => n6504);
   U20982 : OAI22_X1 port map( A1 => n30690, A2 => n26056, B1 => n31041, B2 => 
                           n30682, ZN => n6505);
   U20983 : OAI22_X1 port map( A1 => n30690, A2 => n26055, B1 => n31044, B2 => 
                           n30682, ZN => n6506);
   U20984 : OAI22_X1 port map( A1 => n30690, A2 => n26054, B1 => n31047, B2 => 
                           n30682, ZN => n6507);
   U20985 : OAI22_X1 port map( A1 => n30690, A2 => n26053, B1 => n31050, B2 => 
                           n30682, ZN => n6508);
   U20986 : OAI22_X1 port map( A1 => n30690, A2 => n26052, B1 => n31053, B2 => 
                           n30683, ZN => n6509);
   U20987 : OAI22_X1 port map( A1 => n30690, A2 => n26051, B1 => n31056, B2 => 
                           n30683, ZN => n6510);
   U20988 : OAI22_X1 port map( A1 => n30704, A2 => n25984, B1 => n31059, B2 => 
                           n30696, ZN => n6575);
   U20989 : OAI22_X1 port map( A1 => n30704, A2 => n25983, B1 => n31062, B2 => 
                           n30696, ZN => n6576);
   U20990 : OAI22_X1 port map( A1 => n30704, A2 => n25982, B1 => n31065, B2 => 
                           n30696, ZN => n6577);
   U20991 : OAI22_X1 port map( A1 => n30704, A2 => n25981, B1 => n31068, B2 => 
                           n30696, ZN => n6578);
   U20992 : OAI22_X1 port map( A1 => n30704, A2 => n25980, B1 => n31071, B2 => 
                           n30696, ZN => n6579);
   U20993 : OAI22_X1 port map( A1 => n30704, A2 => n25979, B1 => n31074, B2 => 
                           n30696, ZN => n6580);
   U20994 : OAI22_X1 port map( A1 => n30704, A2 => n25978, B1 => n31077, B2 => 
                           n30696, ZN => n6581);
   U20995 : OAI22_X1 port map( A1 => n30704, A2 => n25977, B1 => n31080, B2 => 
                           n30696, ZN => n6582);
   U20996 : OAI22_X1 port map( A1 => n30704, A2 => n25976, B1 => n31083, B2 => 
                           n30696, ZN => n6583);
   U20997 : OAI22_X1 port map( A1 => n30704, A2 => n25975, B1 => n31086, B2 => 
                           n30696, ZN => n6584);
   U20998 : OAI22_X1 port map( A1 => n30704, A2 => n25974, B1 => n31089, B2 => 
                           n30697, ZN => n6585);
   U20999 : OAI22_X1 port map( A1 => n30704, A2 => n25973, B1 => n31092, B2 => 
                           n30697, ZN => n6586);
   U21000 : OAI22_X1 port map( A1 => n30704, A2 => n25972, B1 => n31095, B2 => 
                           n30697, ZN => n6587);
   U21001 : OAI22_X1 port map( A1 => n30705, A2 => n25971, B1 => n31098, B2 => 
                           n30697, ZN => n6588);
   U21002 : OAI22_X1 port map( A1 => n30705, A2 => n25970, B1 => n31101, B2 => 
                           n30697, ZN => n6589);
   U21003 : OAI22_X1 port map( A1 => n30705, A2 => n25969, B1 => n31104, B2 => 
                           n30697, ZN => n6590);
   U21004 : OAI22_X1 port map( A1 => n30705, A2 => n25968, B1 => n31107, B2 => 
                           n30697, ZN => n6591);
   U21005 : OAI22_X1 port map( A1 => n30705, A2 => n25967, B1 => n31110, B2 => 
                           n30697, ZN => n6592);
   U21006 : OAI22_X1 port map( A1 => n30705, A2 => n25966, B1 => n31113, B2 => 
                           n30697, ZN => n6593);
   U21007 : OAI22_X1 port map( A1 => n30705, A2 => n25965, B1 => n31116, B2 => 
                           n30697, ZN => n6594);
   U21008 : OAI22_X1 port map( A1 => n30705, A2 => n25964, B1 => n31119, B2 => 
                           n30697, ZN => n6595);
   U21009 : OAI22_X1 port map( A1 => n30705, A2 => n25963, B1 => n31122, B2 => 
                           n30697, ZN => n6596);
   U21010 : OAI22_X1 port map( A1 => n30691, A2 => n26050, B1 => n31059, B2 => 
                           n30683, ZN => n6511);
   U21011 : OAI22_X1 port map( A1 => n30691, A2 => n26049, B1 => n31062, B2 => 
                           n30683, ZN => n6512);
   U21012 : OAI22_X1 port map( A1 => n30691, A2 => n26048, B1 => n31065, B2 => 
                           n30683, ZN => n6513);
   U21013 : OAI22_X1 port map( A1 => n30691, A2 => n26047, B1 => n31068, B2 => 
                           n30683, ZN => n6514);
   U21014 : OAI22_X1 port map( A1 => n30691, A2 => n26046, B1 => n31071, B2 => 
                           n30683, ZN => n6515);
   U21015 : OAI22_X1 port map( A1 => n30691, A2 => n26045, B1 => n31074, B2 => 
                           n30683, ZN => n6516);
   U21016 : OAI22_X1 port map( A1 => n30691, A2 => n26044, B1 => n31077, B2 => 
                           n30683, ZN => n6517);
   U21017 : OAI22_X1 port map( A1 => n30691, A2 => n26043, B1 => n31080, B2 => 
                           n30683, ZN => n6518);
   U21018 : OAI22_X1 port map( A1 => n30691, A2 => n26042, B1 => n31083, B2 => 
                           n30683, ZN => n6519);
   U21019 : OAI22_X1 port map( A1 => n30691, A2 => n26041, B1 => n31086, B2 => 
                           n30683, ZN => n6520);
   U21020 : OAI22_X1 port map( A1 => n30691, A2 => n26040, B1 => n31089, B2 => 
                           n30684, ZN => n6521);
   U21021 : OAI22_X1 port map( A1 => n30691, A2 => n26039, B1 => n31092, B2 => 
                           n30684, ZN => n6522);
   U21022 : OAI22_X1 port map( A1 => n30691, A2 => n26038, B1 => n31095, B2 => 
                           n30684, ZN => n6523);
   U21023 : OAI22_X1 port map( A1 => n30692, A2 => n26037, B1 => n31098, B2 => 
                           n30684, ZN => n6524);
   U21024 : OAI22_X1 port map( A1 => n30692, A2 => n26036, B1 => n31101, B2 => 
                           n30684, ZN => n6525);
   U21025 : OAI22_X1 port map( A1 => n30692, A2 => n26035, B1 => n31104, B2 => 
                           n30684, ZN => n6526);
   U21026 : OAI22_X1 port map( A1 => n30692, A2 => n26034, B1 => n31107, B2 => 
                           n30684, ZN => n6527);
   U21027 : OAI22_X1 port map( A1 => n30692, A2 => n26033, B1 => n31110, B2 => 
                           n30684, ZN => n6528);
   U21028 : OAI22_X1 port map( A1 => n30692, A2 => n26032, B1 => n31113, B2 => 
                           n30684, ZN => n6529);
   U21029 : OAI22_X1 port map( A1 => n30692, A2 => n26031, B1 => n31116, B2 => 
                           n30684, ZN => n6530);
   U21030 : OAI22_X1 port map( A1 => n30692, A2 => n26030, B1 => n31119, B2 => 
                           n30684, ZN => n6531);
   U21031 : OAI22_X1 port map( A1 => n30692, A2 => n26029, B1 => n31122, B2 => 
                           n30684, ZN => n6532);
   U21032 : OAI22_X1 port map( A1 => n30565, A2 => n27678, B1 => n30980, B2 => 
                           n30557, ZN => n5794);
   U21033 : OAI22_X1 port map( A1 => n30565, A2 => n27652, B1 => n30983, B2 => 
                           n30557, ZN => n5796);
   U21034 : OAI22_X1 port map( A1 => n30565, A2 => n27626, B1 => n30986, B2 => 
                           n30557, ZN => n5798);
   U21035 : OAI22_X1 port map( A1 => n30565, A2 => n27600, B1 => n30989, B2 => 
                           n30557, ZN => n5800);
   U21036 : OAI22_X1 port map( A1 => n30565, A2 => n27574, B1 => n30992, B2 => 
                           n30557, ZN => n5802);
   U21037 : OAI22_X1 port map( A1 => n30565, A2 => n27548, B1 => n30995, B2 => 
                           n30557, ZN => n5804);
   U21038 : OAI22_X1 port map( A1 => n30565, A2 => n27522, B1 => n30998, B2 => 
                           n30557, ZN => n5806);
   U21039 : OAI22_X1 port map( A1 => n30565, A2 => n27496, B1 => n31001, B2 => 
                           n30557, ZN => n5808);
   U21040 : OAI22_X1 port map( A1 => n30565, A2 => n27470, B1 => n31004, B2 => 
                           n30557, ZN => n5810);
   U21041 : OAI22_X1 port map( A1 => n30565, A2 => n27444, B1 => n31007, B2 => 
                           n30557, ZN => n5812);
   U21042 : OAI22_X1 port map( A1 => n30565, A2 => n27418, B1 => n31010, B2 => 
                           n30557, ZN => n5814);
   U21043 : OAI22_X1 port map( A1 => n30565, A2 => n27392, B1 => n31013, B2 => 
                           n30557, ZN => n5816);
   U21044 : OAI22_X1 port map( A1 => n30565, A2 => n27366, B1 => n31016, B2 => 
                           n30558, ZN => n5818);
   U21045 : OAI22_X1 port map( A1 => n30566, A2 => n27340, B1 => n31019, B2 => 
                           n30558, ZN => n5820);
   U21046 : OAI22_X1 port map( A1 => n30566, A2 => n27314, B1 => n31022, B2 => 
                           n30558, ZN => n5822);
   U21047 : OAI22_X1 port map( A1 => n30566, A2 => n27288, B1 => n31025, B2 => 
                           n30558, ZN => n5824);
   U21048 : OAI22_X1 port map( A1 => n30566, A2 => n27262, B1 => n31028, B2 => 
                           n30558, ZN => n5826);
   U21049 : OAI22_X1 port map( A1 => n30566, A2 => n27236, B1 => n31031, B2 => 
                           n30558, ZN => n5828);
   U21050 : OAI22_X1 port map( A1 => n30566, A2 => n27210, B1 => n31034, B2 => 
                           n30558, ZN => n5830);
   U21051 : OAI22_X1 port map( A1 => n30566, A2 => n27184, B1 => n31037, B2 => 
                           n30558, ZN => n5832);
   U21052 : OAI22_X1 port map( A1 => n30566, A2 => n27158, B1 => n31040, B2 => 
                           n30558, ZN => n5834);
   U21053 : OAI22_X1 port map( A1 => n30566, A2 => n27132, B1 => n31043, B2 => 
                           n30558, ZN => n5836);
   U21054 : OAI22_X1 port map( A1 => n30566, A2 => n27106, B1 => n31046, B2 => 
                           n30558, ZN => n5838);
   U21055 : OAI22_X1 port map( A1 => n30566, A2 => n27080, B1 => n31049, B2 => 
                           n30558, ZN => n5840);
   U21056 : OAI22_X1 port map( A1 => n30566, A2 => n27054, B1 => n31052, B2 => 
                           n30559, ZN => n5842);
   U21057 : OAI22_X1 port map( A1 => n30566, A2 => n27028, B1 => n31055, B2 => 
                           n30559, ZN => n5844);
   U21058 : OAI22_X1 port map( A1 => n30567, A2 => n27002, B1 => n31058, B2 => 
                           n30559, ZN => n5846);
   U21059 : OAI22_X1 port map( A1 => n30567, A2 => n26976, B1 => n31061, B2 => 
                           n30559, ZN => n5848);
   U21060 : OAI22_X1 port map( A1 => n30567, A2 => n26950, B1 => n31064, B2 => 
                           n30559, ZN => n5850);
   U21061 : OAI22_X1 port map( A1 => n30567, A2 => n26924, B1 => n31067, B2 => 
                           n30559, ZN => n5852);
   U21062 : OAI22_X1 port map( A1 => n30567, A2 => n26898, B1 => n31070, B2 => 
                           n30559, ZN => n5854);
   U21063 : OAI22_X1 port map( A1 => n30567, A2 => n26872, B1 => n31073, B2 => 
                           n30559, ZN => n5856);
   U21064 : OAI22_X1 port map( A1 => n30567, A2 => n26846, B1 => n31076, B2 => 
                           n30559, ZN => n5858);
   U21065 : OAI22_X1 port map( A1 => n30567, A2 => n26820, B1 => n31079, B2 => 
                           n30559, ZN => n5860);
   U21066 : OAI22_X1 port map( A1 => n30567, A2 => n26794, B1 => n31082, B2 => 
                           n30559, ZN => n5862);
   U21067 : OAI22_X1 port map( A1 => n30567, A2 => n26768, B1 => n31085, B2 => 
                           n30559, ZN => n5864);
   U21068 : OAI22_X1 port map( A1 => n30567, A2 => n26742, B1 => n31088, B2 => 
                           n30560, ZN => n5866);
   U21069 : OAI22_X1 port map( A1 => n30567, A2 => n26716, B1 => n31091, B2 => 
                           n30560, ZN => n5868);
   U21070 : OAI22_X1 port map( A1 => n30567, A2 => n26690, B1 => n31094, B2 => 
                           n30560, ZN => n5870);
   U21071 : OAI22_X1 port map( A1 => n30568, A2 => n26664, B1 => n31097, B2 => 
                           n30560, ZN => n5872);
   U21072 : OAI22_X1 port map( A1 => n30568, A2 => n26638, B1 => n31100, B2 => 
                           n30560, ZN => n5874);
   U21073 : OAI22_X1 port map( A1 => n30568, A2 => n26612, B1 => n31103, B2 => 
                           n30560, ZN => n5876);
   U21074 : OAI22_X1 port map( A1 => n30568, A2 => n26586, B1 => n31106, B2 => 
                           n30560, ZN => n5878);
   U21075 : OAI22_X1 port map( A1 => n30568, A2 => n26560, B1 => n31109, B2 => 
                           n30560, ZN => n5880);
   U21076 : OAI22_X1 port map( A1 => n30568, A2 => n26534, B1 => n31112, B2 => 
                           n30560, ZN => n5882);
   U21077 : OAI22_X1 port map( A1 => n30568, A2 => n26508, B1 => n31115, B2 => 
                           n30560, ZN => n5884);
   U21078 : OAI22_X1 port map( A1 => n30568, A2 => n26482, B1 => n31118, B2 => 
                           n30560, ZN => n5886);
   U21079 : OAI22_X1 port map( A1 => n30568, A2 => n26456, B1 => n31121, B2 => 
                           n30560, ZN => n5888);
   U21080 : OAI22_X1 port map( A1 => n30701, A2 => n26022, B1 => n30945, B2 => 
                           n30693, ZN => n6537);
   U21081 : OAI22_X1 port map( A1 => n30701, A2 => n26021, B1 => n30948, B2 => 
                           n30693, ZN => n6538);
   U21082 : OAI22_X1 port map( A1 => n30701, A2 => n26020, B1 => n30951, B2 => 
                           n30693, ZN => n6539);
   U21083 : OAI22_X1 port map( A1 => n30701, A2 => n26019, B1 => n30954, B2 => 
                           n30693, ZN => n6540);
   U21084 : OAI22_X1 port map( A1 => n30701, A2 => n26018, B1 => n30957, B2 => 
                           n30693, ZN => n6541);
   U21085 : OAI22_X1 port map( A1 => n30701, A2 => n26017, B1 => n30960, B2 => 
                           n30693, ZN => n6542);
   U21086 : OAI22_X1 port map( A1 => n30701, A2 => n26016, B1 => n30963, B2 => 
                           n30693, ZN => n6543);
   U21087 : OAI22_X1 port map( A1 => n30701, A2 => n26015, B1 => n30966, B2 => 
                           n30693, ZN => n6544);
   U21088 : OAI22_X1 port map( A1 => n30701, A2 => n26014, B1 => n30969, B2 => 
                           n30693, ZN => n6545);
   U21089 : OAI22_X1 port map( A1 => n30701, A2 => n26013, B1 => n30972, B2 => 
                           n30693, ZN => n6546);
   U21090 : OAI22_X1 port map( A1 => n30701, A2 => n26012, B1 => n30975, B2 => 
                           n30693, ZN => n6547);
   U21091 : OAI22_X1 port map( A1 => n30701, A2 => n26011, B1 => n30978, B2 => 
                           n30693, ZN => n6548);
   U21092 : OAI22_X1 port map( A1 => n30688, A2 => n26088, B1 => n30945, B2 => 
                           n30680, ZN => n6473);
   U21093 : OAI22_X1 port map( A1 => n30688, A2 => n26087, B1 => n30948, B2 => 
                           n30680, ZN => n6474);
   U21094 : OAI22_X1 port map( A1 => n30688, A2 => n26086, B1 => n30951, B2 => 
                           n30680, ZN => n6475);
   U21095 : OAI22_X1 port map( A1 => n30688, A2 => n26085, B1 => n30954, B2 => 
                           n30680, ZN => n6476);
   U21096 : OAI22_X1 port map( A1 => n30688, A2 => n26084, B1 => n30957, B2 => 
                           n30680, ZN => n6477);
   U21097 : OAI22_X1 port map( A1 => n30688, A2 => n26083, B1 => n30960, B2 => 
                           n30680, ZN => n6478);
   U21098 : OAI22_X1 port map( A1 => n30688, A2 => n26082, B1 => n30963, B2 => 
                           n30680, ZN => n6479);
   U21099 : OAI22_X1 port map( A1 => n30688, A2 => n26081, B1 => n30966, B2 => 
                           n30680, ZN => n6480);
   U21100 : OAI22_X1 port map( A1 => n30688, A2 => n26080, B1 => n30969, B2 => 
                           n30680, ZN => n6481);
   U21101 : OAI22_X1 port map( A1 => n30688, A2 => n26079, B1 => n30972, B2 => 
                           n30680, ZN => n6482);
   U21102 : OAI22_X1 port map( A1 => n30688, A2 => n26078, B1 => n30975, B2 => 
                           n30680, ZN => n6483);
   U21103 : OAI22_X1 port map( A1 => n30688, A2 => n26077, B1 => n30978, B2 => 
                           n30680, ZN => n6484);
   U21104 : OAI22_X1 port map( A1 => n30564, A2 => n27990, B1 => n30944, B2 => 
                           n30556, ZN => n5770);
   U21105 : OAI22_X1 port map( A1 => n30564, A2 => n27964, B1 => n30947, B2 => 
                           n30556, ZN => n5772);
   U21106 : OAI22_X1 port map( A1 => n30564, A2 => n27938, B1 => n30950, B2 => 
                           n30556, ZN => n5774);
   U21107 : OAI22_X1 port map( A1 => n30564, A2 => n27912, B1 => n30953, B2 => 
                           n30556, ZN => n5776);
   U21108 : OAI22_X1 port map( A1 => n30564, A2 => n27886, B1 => n30956, B2 => 
                           n30556, ZN => n5778);
   U21109 : OAI22_X1 port map( A1 => n30564, A2 => n27860, B1 => n30959, B2 => 
                           n30556, ZN => n5780);
   U21110 : OAI22_X1 port map( A1 => n30564, A2 => n27834, B1 => n30962, B2 => 
                           n30556, ZN => n5782);
   U21111 : OAI22_X1 port map( A1 => n30564, A2 => n27808, B1 => n30965, B2 => 
                           n30556, ZN => n5784);
   U21112 : OAI22_X1 port map( A1 => n30564, A2 => n27782, B1 => n30968, B2 => 
                           n30556, ZN => n5786);
   U21113 : OAI22_X1 port map( A1 => n30564, A2 => n27756, B1 => n30971, B2 => 
                           n30556, ZN => n5788);
   U21114 : OAI22_X1 port map( A1 => n30564, A2 => n27730, B1 => n30974, B2 => 
                           n30556, ZN => n5790);
   U21115 : OAI22_X1 port map( A1 => n30564, A2 => n27704, B1 => n30977, B2 => 
                           n30556, ZN => n5792);
   U21116 : OAI22_X1 port map( A1 => n30728, A2 => n25950, B1 => n30957, B2 => 
                           n30718, ZN => n6669);
   U21117 : OAI22_X1 port map( A1 => n30728, A2 => n25949, B1 => n30960, B2 => 
                           n30718, ZN => n6670);
   U21118 : OAI22_X1 port map( A1 => n30728, A2 => n25948, B1 => n30963, B2 => 
                           n30718, ZN => n6671);
   U21119 : OAI22_X1 port map( A1 => n30728, A2 => n25947, B1 => n30966, B2 => 
                           n30718, ZN => n6672);
   U21120 : OAI22_X1 port map( A1 => n30728, A2 => n25946, B1 => n30969, B2 => 
                           n30718, ZN => n6673);
   U21121 : OAI22_X1 port map( A1 => n30728, A2 => n25945, B1 => n30972, B2 => 
                           n30718, ZN => n6674);
   U21122 : OAI22_X1 port map( A1 => n30728, A2 => n25944, B1 => n30975, B2 => 
                           n30718, ZN => n6675);
   U21123 : OAI22_X1 port map( A1 => n30728, A2 => n25943, B1 => n30978, B2 => 
                           n30718, ZN => n6676);
   U21124 : OAI22_X1 port map( A1 => n30729, A2 => n25954, B1 => n30945, B2 => 
                           n30718, ZN => n6665);
   U21125 : OAI22_X1 port map( A1 => n30729, A2 => n25953, B1 => n30948, B2 => 
                           n30718, ZN => n6666);
   U21126 : OAI22_X1 port map( A1 => n30729, A2 => n25952, B1 => n30951, B2 => 
                           n30718, ZN => n6667);
   U21127 : OAI22_X1 port map( A1 => n30729, A2 => n25951, B1 => n30954, B2 => 
                           n30718, ZN => n6668);
   U21128 : OAI22_X1 port map( A1 => n30788, A2 => n25801, B1 => n30945, B2 => 
                           n30780, ZN => n6985);
   U21129 : OAI22_X1 port map( A1 => n30788, A2 => n25800, B1 => n30948, B2 => 
                           n30780, ZN => n6986);
   U21130 : OAI22_X1 port map( A1 => n30788, A2 => n25799, B1 => n30951, B2 => 
                           n30780, ZN => n6987);
   U21131 : OAI22_X1 port map( A1 => n30788, A2 => n25798, B1 => n30954, B2 => 
                           n30780, ZN => n6988);
   U21132 : OAI22_X1 port map( A1 => n30788, A2 => n25797, B1 => n30957, B2 => 
                           n30780, ZN => n6989);
   U21133 : OAI22_X1 port map( A1 => n30788, A2 => n25796, B1 => n30960, B2 => 
                           n30780, ZN => n6990);
   U21134 : OAI22_X1 port map( A1 => n30788, A2 => n25795, B1 => n30963, B2 => 
                           n30780, ZN => n6991);
   U21135 : OAI22_X1 port map( A1 => n30788, A2 => n25794, B1 => n30966, B2 => 
                           n30780, ZN => n6992);
   U21136 : OAI22_X1 port map( A1 => n30788, A2 => n25793, B1 => n30969, B2 => 
                           n30780, ZN => n6993);
   U21137 : OAI22_X1 port map( A1 => n30788, A2 => n25792, B1 => n30972, B2 => 
                           n30780, ZN => n6994);
   U21138 : OAI22_X1 port map( A1 => n30788, A2 => n25791, B1 => n30975, B2 => 
                           n30780, ZN => n6995);
   U21139 : OAI22_X1 port map( A1 => n30788, A2 => n25790, B1 => n30978, B2 => 
                           n30780, ZN => n6996);
   U21140 : OAI22_X1 port map( A1 => n30789, A2 => n25789, B1 => n30981, B2 => 
                           n30781, ZN => n6997);
   U21141 : OAI22_X1 port map( A1 => n30789, A2 => n25788, B1 => n30984, B2 => 
                           n30781, ZN => n6998);
   U21142 : OAI22_X1 port map( A1 => n30789, A2 => n25787, B1 => n30987, B2 => 
                           n30781, ZN => n6999);
   U21143 : OAI22_X1 port map( A1 => n30789, A2 => n25786, B1 => n30990, B2 => 
                           n30781, ZN => n7000);
   U21144 : OAI22_X1 port map( A1 => n30789, A2 => n25785, B1 => n30993, B2 => 
                           n30781, ZN => n7001);
   U21145 : OAI22_X1 port map( A1 => n30789, A2 => n25784, B1 => n30996, B2 => 
                           n30781, ZN => n7002);
   U21146 : OAI22_X1 port map( A1 => n30789, A2 => n25783, B1 => n30999, B2 => 
                           n30781, ZN => n7003);
   U21147 : OAI22_X1 port map( A1 => n30789, A2 => n25782, B1 => n31002, B2 => 
                           n30781, ZN => n7004);
   U21148 : OAI22_X1 port map( A1 => n30789, A2 => n25781, B1 => n31005, B2 => 
                           n30781, ZN => n7005);
   U21149 : OAI22_X1 port map( A1 => n30789, A2 => n25780, B1 => n31008, B2 => 
                           n30781, ZN => n7006);
   U21150 : OAI22_X1 port map( A1 => n30789, A2 => n25779, B1 => n31011, B2 => 
                           n30781, ZN => n7007);
   U21151 : OAI22_X1 port map( A1 => n30789, A2 => n25778, B1 => n31014, B2 => 
                           n30781, ZN => n7008);
   U21152 : OAI22_X1 port map( A1 => n30789, A2 => n25777, B1 => n31017, B2 => 
                           n30782, ZN => n7009);
   U21153 : OAI22_X1 port map( A1 => n30790, A2 => n25776, B1 => n31020, B2 => 
                           n30782, ZN => n7010);
   U21154 : OAI22_X1 port map( A1 => n30790, A2 => n25775, B1 => n31023, B2 => 
                           n30782, ZN => n7011);
   U21155 : OAI22_X1 port map( A1 => n30790, A2 => n25774, B1 => n31026, B2 => 
                           n30782, ZN => n7012);
   U21156 : OAI22_X1 port map( A1 => n30790, A2 => n25773, B1 => n31029, B2 => 
                           n30782, ZN => n7013);
   U21157 : OAI22_X1 port map( A1 => n30790, A2 => n25772, B1 => n31032, B2 => 
                           n30782, ZN => n7014);
   U21158 : OAI22_X1 port map( A1 => n30790, A2 => n25771, B1 => n31035, B2 => 
                           n30782, ZN => n7015);
   U21159 : OAI22_X1 port map( A1 => n30790, A2 => n25770, B1 => n31038, B2 => 
                           n30782, ZN => n7016);
   U21160 : OAI22_X1 port map( A1 => n30790, A2 => n25769, B1 => n31041, B2 => 
                           n30782, ZN => n7017);
   U21161 : OAI22_X1 port map( A1 => n30790, A2 => n25768, B1 => n31044, B2 => 
                           n30782, ZN => n7018);
   U21162 : OAI22_X1 port map( A1 => n30790, A2 => n25767, B1 => n31047, B2 => 
                           n30782, ZN => n7019);
   U21163 : OAI22_X1 port map( A1 => n30790, A2 => n25766, B1 => n31050, B2 => 
                           n30782, ZN => n7020);
   U21164 : OAI22_X1 port map( A1 => n30790, A2 => n25765, B1 => n31053, B2 => 
                           n30783, ZN => n7021);
   U21165 : OAI22_X1 port map( A1 => n30790, A2 => n25764, B1 => n31056, B2 => 
                           n30783, ZN => n7022);
   U21166 : OAI22_X1 port map( A1 => n30791, A2 => n25763, B1 => n31059, B2 => 
                           n30783, ZN => n7023);
   U21167 : OAI22_X1 port map( A1 => n30791, A2 => n25762, B1 => n31062, B2 => 
                           n30783, ZN => n7024);
   U21168 : OAI22_X1 port map( A1 => n30791, A2 => n25761, B1 => n31065, B2 => 
                           n30783, ZN => n7025);
   U21169 : OAI22_X1 port map( A1 => n30791, A2 => n25760, B1 => n31068, B2 => 
                           n30783, ZN => n7026);
   U21170 : OAI22_X1 port map( A1 => n30791, A2 => n25759, B1 => n31071, B2 => 
                           n30783, ZN => n7027);
   U21171 : OAI22_X1 port map( A1 => n30791, A2 => n25758, B1 => n31074, B2 => 
                           n30783, ZN => n7028);
   U21172 : OAI22_X1 port map( A1 => n30791, A2 => n25757, B1 => n31077, B2 => 
                           n30783, ZN => n7029);
   U21173 : OAI22_X1 port map( A1 => n30791, A2 => n25756, B1 => n31080, B2 => 
                           n30783, ZN => n7030);
   U21174 : OAI22_X1 port map( A1 => n30791, A2 => n25755, B1 => n31083, B2 => 
                           n30783, ZN => n7031);
   U21175 : OAI22_X1 port map( A1 => n30791, A2 => n25754, B1 => n31086, B2 => 
                           n30783, ZN => n7032);
   U21176 : OAI22_X1 port map( A1 => n30791, A2 => n25753, B1 => n31089, B2 => 
                           n30784, ZN => n7033);
   U21177 : OAI22_X1 port map( A1 => n30791, A2 => n25752, B1 => n31092, B2 => 
                           n30784, ZN => n7034);
   U21178 : OAI22_X1 port map( A1 => n30791, A2 => n25751, B1 => n31095, B2 => 
                           n30784, ZN => n7035);
   U21179 : OAI22_X1 port map( A1 => n30792, A2 => n25750, B1 => n31098, B2 => 
                           n30784, ZN => n7036);
   U21180 : OAI22_X1 port map( A1 => n30792, A2 => n25749, B1 => n31101, B2 => 
                           n30784, ZN => n7037);
   U21181 : OAI22_X1 port map( A1 => n30792, A2 => n25748, B1 => n31104, B2 => 
                           n30784, ZN => n7038);
   U21182 : OAI22_X1 port map( A1 => n30792, A2 => n25747, B1 => n31107, B2 => 
                           n30784, ZN => n7039);
   U21183 : OAI22_X1 port map( A1 => n30792, A2 => n25746, B1 => n31110, B2 => 
                           n30784, ZN => n7040);
   U21184 : OAI22_X1 port map( A1 => n30792, A2 => n25745, B1 => n31113, B2 => 
                           n30784, ZN => n7041);
   U21185 : OAI22_X1 port map( A1 => n30792, A2 => n25744, B1 => n31116, B2 => 
                           n30784, ZN => n7042);
   U21186 : OAI22_X1 port map( A1 => n30792, A2 => n25743, B1 => n31119, B2 => 
                           n30784, ZN => n7043);
   U21187 : OAI22_X1 port map( A1 => n30792, A2 => n25742, B1 => n31122, B2 => 
                           n30784, ZN => n7044);
   U21188 : OAI21_X1 port map( B1 => n25235, B2 => n25451, A => n31163, ZN => 
                           n25455);
   U21189 : OAI21_X1 port map( B1 => n25235, B2 => n25302, A => n31163, ZN => 
                           n25303);
   U21190 : OAI21_X1 port map( B1 => n25231, B2 => n25302, A => n31163, ZN => 
                           n25236);
   U21191 : OAI21_X1 port map( B1 => n25231, B2 => n25451, A => n31163, ZN => 
                           n25385);
   U21192 : OAI21_X1 port map( B1 => n25232, B2 => n25587, A => n31163, ZN => 
                           n25521);
   U21193 : OAI21_X1 port map( B1 => n25382, B2 => n25587, A => n31163, ZN => 
                           n25670);
   U21194 : OAI21_X1 port map( B1 => n25382, B2 => n25654, A => n31161, ZN => 
                           n25736);
   U21195 : OAI21_X1 port map( B1 => n25232, B2 => n25654, A => n31162, ZN => 
                           n25588);
   U21196 : OAI21_X1 port map( B1 => n25451, B2 => n26099, A => n31161, ZN => 
                           n26316);
   U21197 : OAI21_X1 port map( B1 => n25382, B2 => n25873, A => n31162, ZN => 
                           n25957);
   U21198 : OAI21_X1 port map( B1 => n25302, B2 => n26099, A => n31161, ZN => 
                           n26168);
   U21199 : OAI21_X1 port map( B1 => n25382, B2 => n25940, A => n31161, ZN => 
                           n26023);
   U21200 : OAI21_X1 port map( B1 => n25302, B2 => n26096, A => n31161, ZN => 
                           n26102);
   U21201 : OAI21_X1 port map( B1 => n25451, B2 => n26096, A => n31161, ZN => 
                           n26250);
   U21202 : OAI21_X1 port map( B1 => n25232, B2 => n25940, A => n31161, ZN => 
                           n25874);
   U21203 : AND2_X1 port map( A1 => n29284, A2 => n29300, ZN => n28073);
   U21204 : AND2_X1 port map( A1 => n29284, A2 => n29299, ZN => n28074);
   U21205 : AND2_X1 port map( A1 => n28001, A2 => n28020, ZN => n26352);
   U21206 : AND2_X1 port map( A1 => n28001, A2 => n28019, ZN => n26353);
   U21207 : AND2_X1 port map( A1 => n29282, A2 => n29303, ZN => n28078);
   U21208 : AND2_X1 port map( A1 => n29282, A2 => n29302, ZN => n28079);
   U21209 : AND2_X1 port map( A1 => n29282, A2 => n29300, ZN => n28083);
   U21210 : AND2_X1 port map( A1 => n29282, A2 => n29299, ZN => n28084);
   U21211 : AND2_X1 port map( A1 => n29302, A2 => n29287, ZN => n28089);
   U21212 : AND2_X1 port map( A1 => n28009, A2 => n28001, ZN => n26339);
   U21213 : AND2_X1 port map( A1 => n28006, A2 => n28020, ZN => n26371);
   U21214 : AND2_X1 port map( A1 => n28006, A2 => n28019, ZN => n26373);
   U21215 : AND2_X1 port map( A1 => n28006, A2 => n28010, ZN => n26357);
   U21216 : AND2_X1 port map( A1 => n28006, A2 => n28009, ZN => n26359);
   U21217 : AND2_X1 port map( A1 => n29303, A2 => n29287, ZN => n28088);
   U21218 : AND2_X1 port map( A1 => n28010, A2 => n28001, ZN => n26338);
   U21219 : AND2_X1 port map( A1 => n29283, A2 => n29287, ZN => n28054);
   U21220 : AND2_X1 port map( A1 => n29281, A2 => n29287, ZN => n28055);
   U21221 : AND2_X1 port map( A1 => n29283, A2 => n29284, ZN => n28049);
   U21222 : AND2_X1 port map( A1 => n29281, A2 => n29284, ZN => n28050);
   U21223 : AND2_X1 port map( A1 => n29291, A2 => n29286, ZN => n28059);
   U21224 : AND2_X1 port map( A1 => n29290, A2 => n29286, ZN => n28060);
   U21225 : AND2_X1 port map( A1 => n29291, A2 => n29282, ZN => n28064);
   U21226 : AND2_X1 port map( A1 => n29290, A2 => n29282, ZN => n28065);
   U21227 : AND2_X1 port map( A1 => n28013, A2 => n28003, ZN => n26343);
   U21228 : AND2_X1 port map( A1 => n28012, A2 => n28003, ZN => n26344);
   U21229 : AND2_X1 port map( A1 => n28002, A2 => n28006, ZN => n26333);
   U21230 : AND2_X1 port map( A1 => n28000, A2 => n28006, ZN => n26334);
   U21231 : AND2_X1 port map( A1 => n28002, A2 => n28003, ZN => n26328);
   U21232 : AND2_X1 port map( A1 => n28000, A2 => n28003, ZN => n26329);
   U21233 : AND2_X1 port map( A1 => n28013, A2 => n28001, ZN => n26364);
   U21234 : AND2_X1 port map( A1 => n28012, A2 => n28001, ZN => n26366);
   U21235 : AND2_X1 port map( A1 => n29275, A2 => n31187, ZN => n28044);
   U21236 : AND2_X1 port map( A1 => n27994, A2 => n31187, ZN => n26323);
   U21237 : BUF_X1 port map( A => n25150, Z => n31159);
   U21238 : BUF_X1 port map( A => n25150, Z => n31160);
   U21239 : NOR2_X1 port map( A1 => n29308, A2 => ADD_RD1(2), ZN => n29284);
   U21240 : NOR2_X1 port map( A1 => n28033, A2 => ADD_RD2(2), ZN => n28003);
   U21241 : NOR3_X1 port map( A1 => n29306, A2 => ADD_RD1(0), A3 => n29293, ZN 
                           => n29299);
   U21242 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(3), A3 => n28029,
                           ZN => n28019);
   U21243 : NOR2_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), ZN => n28001)
                           ;
   U21244 : NOR3_X1 port map( A1 => n28029, A2 => ADD_RD2(3), A3 => n28007, ZN 
                           => n28020);
   U21245 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(3), A3 => n29306,
                           ZN => n29302);
   U21246 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(4), A3 => n28024,
                           ZN => n28009);
   U21247 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n29282)
                           ;
   U21248 : NOR3_X1 port map( A1 => n28024, A2 => ADD_RD2(4), A3 => n28007, ZN 
                           => n28010);
   U21249 : NOR3_X1 port map( A1 => n29306, A2 => ADD_RD1(3), A3 => n29288, ZN 
                           => n29303);
   U21250 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => 
                           ADD_RD1(0), ZN => n29281);
   U21251 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => 
                           ADD_RD2(0), ZN => n28000);
   U21252 : NOR3_X1 port map( A1 => n29288, A2 => ADD_RD1(4), A3 => n29293, ZN 
                           => n29291);
   U21253 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => n29288,
                           ZN => n29283);
   U21254 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(4), A3 => n29293,
                           ZN => n29290);
   U21255 : NOR3_X1 port map( A1 => n28029, A2 => ADD_RD2(0), A3 => n28024, ZN 
                           => n28012);
   U21256 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => n28007,
                           ZN => n28002);
   U21257 : NOR4_X1 port map( A1 => n25806, A2 => n29313, A3 => n29314, A4 => 
                           n29315, ZN => n29312);
   U21258 : XNOR2_X1 port map( A => n26101, B => ADD_RD1(1), ZN => n29315);
   U21259 : XNOR2_X1 port map( A => ADD_WR(4), B => n29306, ZN => n29314);
   U21260 : NOR4_X1 port map( A1 => n25153, A2 => n25806, A3 => n28038, A4 => 
                           n28039, ZN => n28037);
   U21261 : XNOR2_X1 port map( A => n26101, B => ADD_RD2(1), ZN => n28039);
   U21262 : XNOR2_X1 port map( A => ADD_WR(4), B => n28029, ZN => n28038);
   U21263 : AOI221_X1 port map( B1 => n30237, B2 => n21987, C1 => n30231, C2 =>
                           n9607, A => n29298, ZN => n29297);
   U21264 : OAI22_X1 port map( A1 => n27990, A2 => n30225, B1 => n26315, B2 => 
                           n30219, ZN => n29298);
   U21265 : AOI221_X1 port map( B1 => n30237, B2 => n21988, C1 => n30231, C2 =>
                           n9602, A => n29268, ZN => n29267);
   U21266 : OAI22_X1 port map( A1 => n27964, A2 => n30225, B1 => n26314, B2 => 
                           n30219, ZN => n29268);
   U21267 : AOI221_X1 port map( B1 => n30237, B2 => n21989, C1 => n30231, C2 =>
                           n9597, A => n29249, ZN => n29248);
   U21268 : OAI22_X1 port map( A1 => n27938, A2 => n30225, B1 => n26313, B2 => 
                           n30219, ZN => n29249);
   U21269 : AOI221_X1 port map( B1 => n30237, B2 => n21990, C1 => n30231, C2 =>
                           n9592, A => n29230, ZN => n29229);
   U21270 : OAI22_X1 port map( A1 => n27912, A2 => n30225, B1 => n26312, B2 => 
                           n30219, ZN => n29230);
   U21271 : AOI221_X1 port map( B1 => n30237, B2 => n21991, C1 => n30231, C2 =>
                           n9587, A => n29211, ZN => n29210);
   U21272 : OAI22_X1 port map( A1 => n27886, A2 => n30225, B1 => n26311, B2 => 
                           n30219, ZN => n29211);
   U21273 : AOI221_X1 port map( B1 => n30237, B2 => n21992, C1 => n30231, C2 =>
                           n9582, A => n29192, ZN => n29191);
   U21274 : OAI22_X1 port map( A1 => n27860, A2 => n30225, B1 => n26310, B2 => 
                           n30219, ZN => n29192);
   U21275 : AOI221_X1 port map( B1 => n30237, B2 => n21993, C1 => n30231, C2 =>
                           n9577, A => n29173, ZN => n29172);
   U21276 : OAI22_X1 port map( A1 => n27834, A2 => n30225, B1 => n26309, B2 => 
                           n30219, ZN => n29173);
   U21277 : AOI221_X1 port map( B1 => n30237, B2 => n21994, C1 => n30231, C2 =>
                           n9572, A => n29154, ZN => n29153);
   U21278 : OAI22_X1 port map( A1 => n27808, A2 => n30225, B1 => n26308, B2 => 
                           n30219, ZN => n29154);
   U21279 : AOI221_X1 port map( B1 => n30237, B2 => n21995, C1 => n30231, C2 =>
                           n9567, A => n29135, ZN => n29134);
   U21280 : OAI22_X1 port map( A1 => n27782, A2 => n30225, B1 => n26307, B2 => 
                           n30219, ZN => n29135);
   U21281 : AOI221_X1 port map( B1 => n30237, B2 => n21996, C1 => n30231, C2 =>
                           n9562, A => n29116, ZN => n29115);
   U21282 : OAI22_X1 port map( A1 => n27756, A2 => n30225, B1 => n26306, B2 => 
                           n30219, ZN => n29116);
   U21283 : AOI221_X1 port map( B1 => n30237, B2 => n21997, C1 => n30231, C2 =>
                           n9557, A => n29097, ZN => n29096);
   U21284 : OAI22_X1 port map( A1 => n27730, A2 => n30225, B1 => n26305, B2 => 
                           n30219, ZN => n29097);
   U21285 : AOI221_X1 port map( B1 => n30237, B2 => n21998, C1 => n30231, C2 =>
                           n9552, A => n29078, ZN => n29077);
   U21286 : OAI22_X1 port map( A1 => n27704, A2 => n30225, B1 => n26304, B2 => 
                           n30219, ZN => n29078);
   U21287 : AOI221_X1 port map( B1 => n30238, B2 => n22076, C1 => n30232, C2 =>
                           n9547, A => n29059, ZN => n29058);
   U21288 : OAI22_X1 port map( A1 => n27678, A2 => n30226, B1 => n26303, B2 => 
                           n30220, ZN => n29059);
   U21289 : AOI221_X1 port map( B1 => n30238, B2 => n22077, C1 => n30232, C2 =>
                           n9542, A => n29040, ZN => n29039);
   U21290 : OAI22_X1 port map( A1 => n27652, A2 => n30226, B1 => n26302, B2 => 
                           n30220, ZN => n29040);
   U21291 : AOI221_X1 port map( B1 => n30238, B2 => n22078, C1 => n30232, C2 =>
                           n9537, A => n29021, ZN => n29020);
   U21292 : OAI22_X1 port map( A1 => n27626, A2 => n30226, B1 => n26301, B2 => 
                           n30220, ZN => n29021);
   U21293 : AOI221_X1 port map( B1 => n30238, B2 => n22079, C1 => n30232, C2 =>
                           n9532, A => n29002, ZN => n29001);
   U21294 : OAI22_X1 port map( A1 => n27600, A2 => n30226, B1 => n26300, B2 => 
                           n30220, ZN => n29002);
   U21295 : AOI221_X1 port map( B1 => n30238, B2 => n22080, C1 => n30232, C2 =>
                           n9527, A => n28983, ZN => n28982);
   U21296 : OAI22_X1 port map( A1 => n27574, A2 => n30226, B1 => n26299, B2 => 
                           n30220, ZN => n28983);
   U21297 : AOI221_X1 port map( B1 => n30238, B2 => n22081, C1 => n30232, C2 =>
                           n9522, A => n28964, ZN => n28963);
   U21298 : OAI22_X1 port map( A1 => n27548, A2 => n30226, B1 => n26298, B2 => 
                           n30220, ZN => n28964);
   U21299 : AOI221_X1 port map( B1 => n30238, B2 => n22082, C1 => n30232, C2 =>
                           n9517, A => n28945, ZN => n28944);
   U21300 : OAI22_X1 port map( A1 => n27522, A2 => n30226, B1 => n26297, B2 => 
                           n30220, ZN => n28945);
   U21301 : AOI221_X1 port map( B1 => n30238, B2 => n22083, C1 => n30232, C2 =>
                           n9512, A => n28926, ZN => n28925);
   U21302 : OAI22_X1 port map( A1 => n27496, A2 => n30226, B1 => n26296, B2 => 
                           n30220, ZN => n28926);
   U21303 : AOI221_X1 port map( B1 => n30238, B2 => n22084, C1 => n30232, C2 =>
                           n9507, A => n28907, ZN => n28906);
   U21304 : OAI22_X1 port map( A1 => n27470, A2 => n30226, B1 => n26295, B2 => 
                           n30220, ZN => n28907);
   U21305 : AOI221_X1 port map( B1 => n30238, B2 => n22085, C1 => n30232, C2 =>
                           n9502, A => n28888, ZN => n28887);
   U21306 : OAI22_X1 port map( A1 => n27444, A2 => n30226, B1 => n26294, B2 => 
                           n30220, ZN => n28888);
   U21307 : AOI221_X1 port map( B1 => n30238, B2 => n22086, C1 => n30232, C2 =>
                           n9497, A => n28869, ZN => n28868);
   U21308 : OAI22_X1 port map( A1 => n27418, A2 => n30226, B1 => n26293, B2 => 
                           n30220, ZN => n28869);
   U21309 : AOI221_X1 port map( B1 => n30238, B2 => n22087, C1 => n30232, C2 =>
                           n9492, A => n28850, ZN => n28849);
   U21310 : OAI22_X1 port map( A1 => n27392, A2 => n30226, B1 => n26292, B2 => 
                           n30220, ZN => n28850);
   U21311 : AOI221_X1 port map( B1 => n30239, B2 => n22088, C1 => n30233, C2 =>
                           n9487, A => n28831, ZN => n28830);
   U21312 : OAI22_X1 port map( A1 => n27366, A2 => n30227, B1 => n26291, B2 => 
                           n30221, ZN => n28831);
   U21313 : AOI221_X1 port map( B1 => n30239, B2 => n22089, C1 => n30233, C2 =>
                           n9482, A => n28812, ZN => n28811);
   U21314 : OAI22_X1 port map( A1 => n27340, A2 => n30227, B1 => n26290, B2 => 
                           n30221, ZN => n28812);
   U21315 : AOI221_X1 port map( B1 => n30239, B2 => n22090, C1 => n30233, C2 =>
                           n9477, A => n28793, ZN => n28792);
   U21316 : OAI22_X1 port map( A1 => n27314, A2 => n30227, B1 => n26289, B2 => 
                           n30221, ZN => n28793);
   U21317 : AOI221_X1 port map( B1 => n30239, B2 => n22091, C1 => n30233, C2 =>
                           n9472, A => n28774, ZN => n28773);
   U21318 : OAI22_X1 port map( A1 => n27288, A2 => n30227, B1 => n26288, B2 => 
                           n30221, ZN => n28774);
   U21319 : AOI221_X1 port map( B1 => n30239, B2 => n22092, C1 => n30233, C2 =>
                           n9467, A => n28755, ZN => n28754);
   U21320 : OAI22_X1 port map( A1 => n27262, A2 => n30227, B1 => n26287, B2 => 
                           n30221, ZN => n28755);
   U21321 : AOI221_X1 port map( B1 => n30239, B2 => n22093, C1 => n30233, C2 =>
                           n9462, A => n28736, ZN => n28735);
   U21322 : OAI22_X1 port map( A1 => n27236, A2 => n30227, B1 => n26286, B2 => 
                           n30221, ZN => n28736);
   U21323 : AOI221_X1 port map( B1 => n30239, B2 => n22094, C1 => n30233, C2 =>
                           n9457, A => n28717, ZN => n28716);
   U21324 : OAI22_X1 port map( A1 => n27210, A2 => n30227, B1 => n26285, B2 => 
                           n30221, ZN => n28717);
   U21325 : AOI221_X1 port map( B1 => n30239, B2 => n22095, C1 => n30233, C2 =>
                           n9452, A => n28698, ZN => n28697);
   U21326 : OAI22_X1 port map( A1 => n27184, A2 => n30227, B1 => n26284, B2 => 
                           n30221, ZN => n28698);
   U21327 : AOI221_X1 port map( B1 => n30239, B2 => n22096, C1 => n30233, C2 =>
                           n9447, A => n28679, ZN => n28678);
   U21328 : OAI22_X1 port map( A1 => n27158, A2 => n30227, B1 => n26283, B2 => 
                           n30221, ZN => n28679);
   U21329 : AOI221_X1 port map( B1 => n30239, B2 => n22097, C1 => n30233, C2 =>
                           n9442, A => n28660, ZN => n28659);
   U21330 : OAI22_X1 port map( A1 => n27132, A2 => n30227, B1 => n26282, B2 => 
                           n30221, ZN => n28660);
   U21331 : AOI221_X1 port map( B1 => n30239, B2 => n22098, C1 => n30233, C2 =>
                           n9437, A => n28641, ZN => n28640);
   U21332 : OAI22_X1 port map( A1 => n27106, A2 => n30227, B1 => n26281, B2 => 
                           n30221, ZN => n28641);
   U21333 : AOI221_X1 port map( B1 => n30239, B2 => n22099, C1 => n30233, C2 =>
                           n9432, A => n28622, ZN => n28621);
   U21334 : OAI22_X1 port map( A1 => n27080, A2 => n30227, B1 => n26280, B2 => 
                           n30221, ZN => n28622);
   U21335 : AOI221_X1 port map( B1 => n30240, B2 => n22100, C1 => n30234, C2 =>
                           n9427, A => n28603, ZN => n28602);
   U21336 : OAI22_X1 port map( A1 => n27054, A2 => n30228, B1 => n26279, B2 => 
                           n30222, ZN => n28603);
   U21337 : AOI221_X1 port map( B1 => n30240, B2 => n22101, C1 => n30234, C2 =>
                           n9422, A => n28584, ZN => n28583);
   U21338 : OAI22_X1 port map( A1 => n27028, A2 => n30228, B1 => n26278, B2 => 
                           n30222, ZN => n28584);
   U21339 : AOI221_X1 port map( B1 => n30240, B2 => n22102, C1 => n30234, C2 =>
                           n9417, A => n28565, ZN => n28564);
   U21340 : OAI22_X1 port map( A1 => n27002, A2 => n30228, B1 => n26277, B2 => 
                           n30222, ZN => n28565);
   U21341 : AOI221_X1 port map( B1 => n30240, B2 => n22103, C1 => n30234, C2 =>
                           n9412, A => n28546, ZN => n28545);
   U21342 : OAI22_X1 port map( A1 => n26976, A2 => n30228, B1 => n26276, B2 => 
                           n30222, ZN => n28546);
   U21343 : AOI221_X1 port map( B1 => n30240, B2 => n22104, C1 => n30234, C2 =>
                           n9407, A => n28527, ZN => n28526);
   U21344 : OAI22_X1 port map( A1 => n26950, A2 => n30228, B1 => n26275, B2 => 
                           n30222, ZN => n28527);
   U21345 : AOI221_X1 port map( B1 => n30240, B2 => n22105, C1 => n30234, C2 =>
                           n9402, A => n28508, ZN => n28507);
   U21346 : OAI22_X1 port map( A1 => n26924, A2 => n30228, B1 => n26274, B2 => 
                           n30222, ZN => n28508);
   U21347 : AOI221_X1 port map( B1 => n30240, B2 => n22106, C1 => n30234, C2 =>
                           n9397, A => n28489, ZN => n28488);
   U21348 : OAI22_X1 port map( A1 => n26898, A2 => n30228, B1 => n26273, B2 => 
                           n30222, ZN => n28489);
   U21349 : AOI221_X1 port map( B1 => n30240, B2 => n22107, C1 => n30234, C2 =>
                           n9392, A => n28470, ZN => n28469);
   U21350 : OAI22_X1 port map( A1 => n26872, A2 => n30228, B1 => n26272, B2 => 
                           n30222, ZN => n28470);
   U21351 : AOI221_X1 port map( B1 => n30240, B2 => n22108, C1 => n30234, C2 =>
                           n9387, A => n28451, ZN => n28450);
   U21352 : OAI22_X1 port map( A1 => n26846, A2 => n30228, B1 => n26271, B2 => 
                           n30222, ZN => n28451);
   U21353 : AOI221_X1 port map( B1 => n30240, B2 => n22109, C1 => n30234, C2 =>
                           n9382, A => n28432, ZN => n28431);
   U21354 : OAI22_X1 port map( A1 => n26820, A2 => n30228, B1 => n26270, B2 => 
                           n30222, ZN => n28432);
   U21355 : AOI221_X1 port map( B1 => n30240, B2 => n22110, C1 => n30234, C2 =>
                           n9377, A => n28413, ZN => n28412);
   U21356 : OAI22_X1 port map( A1 => n26794, A2 => n30228, B1 => n26269, B2 => 
                           n30222, ZN => n28413);
   U21357 : AOI221_X1 port map( B1 => n30240, B2 => n22111, C1 => n30234, C2 =>
                           n9372, A => n28394, ZN => n28393);
   U21358 : OAI22_X1 port map( A1 => n26768, A2 => n30228, B1 => n26268, B2 => 
                           n30222, ZN => n28394);
   U21359 : AOI221_X1 port map( B1 => n30241, B2 => n22112, C1 => n30235, C2 =>
                           n9367, A => n28375, ZN => n28374);
   U21360 : OAI22_X1 port map( A1 => n26742, A2 => n30229, B1 => n26267, B2 => 
                           n30223, ZN => n28375);
   U21361 : AOI221_X1 port map( B1 => n30241, B2 => n22113, C1 => n30235, C2 =>
                           n9362, A => n28356, ZN => n28355);
   U21362 : OAI22_X1 port map( A1 => n26716, A2 => n30229, B1 => n26266, B2 => 
                           n30223, ZN => n28356);
   U21363 : AOI221_X1 port map( B1 => n30241, B2 => n22114, C1 => n30235, C2 =>
                           n9357, A => n28337, ZN => n28336);
   U21364 : OAI22_X1 port map( A1 => n26690, A2 => n30229, B1 => n26265, B2 => 
                           n30223, ZN => n28337);
   U21365 : AOI221_X1 port map( B1 => n30241, B2 => n21999, C1 => n30235, C2 =>
                           n9352, A => n28318, ZN => n28317);
   U21366 : OAI22_X1 port map( A1 => n26664, A2 => n30229, B1 => n26264, B2 => 
                           n30223, ZN => n28318);
   U21367 : AOI221_X1 port map( B1 => n30241, B2 => n22000, C1 => n30235, C2 =>
                           n9347, A => n28299, ZN => n28298);
   U21368 : OAI22_X1 port map( A1 => n26638, A2 => n30229, B1 => n26263, B2 => 
                           n30223, ZN => n28299);
   U21369 : AOI221_X1 port map( B1 => n30241, B2 => n22001, C1 => n30235, C2 =>
                           n9342, A => n28280, ZN => n28279);
   U21370 : OAI22_X1 port map( A1 => n26612, A2 => n30229, B1 => n26262, B2 => 
                           n30223, ZN => n28280);
   U21371 : AOI221_X1 port map( B1 => n30241, B2 => n22002, C1 => n30235, C2 =>
                           n9337, A => n28261, ZN => n28260);
   U21372 : OAI22_X1 port map( A1 => n26586, A2 => n30229, B1 => n26261, B2 => 
                           n30223, ZN => n28261);
   U21373 : AOI221_X1 port map( B1 => n30241, B2 => n22003, C1 => n30235, C2 =>
                           n9332, A => n28242, ZN => n28241);
   U21374 : OAI22_X1 port map( A1 => n26560, A2 => n30229, B1 => n26260, B2 => 
                           n30223, ZN => n28242);
   U21375 : AOI221_X1 port map( B1 => n30241, B2 => n22004, C1 => n30235, C2 =>
                           n9327, A => n28223, ZN => n28222);
   U21376 : OAI22_X1 port map( A1 => n26534, A2 => n30229, B1 => n26259, B2 => 
                           n30223, ZN => n28223);
   U21377 : AOI221_X1 port map( B1 => n30241, B2 => n22005, C1 => n30235, C2 =>
                           n9322, A => n28204, ZN => n28203);
   U21378 : OAI22_X1 port map( A1 => n26508, A2 => n30229, B1 => n26258, B2 => 
                           n30223, ZN => n28204);
   U21379 : AOI221_X1 port map( B1 => n30241, B2 => n22006, C1 => n30235, C2 =>
                           n9317, A => n28185, ZN => n28184);
   U21380 : OAI22_X1 port map( A1 => n26482, A2 => n30229, B1 => n26257, B2 => 
                           n30223, ZN => n28185);
   U21381 : AOI221_X1 port map( B1 => n30241, B2 => n22007, C1 => n30235, C2 =>
                           n9312, A => n28166, ZN => n28165);
   U21382 : OAI22_X1 port map( A1 => n26456, A2 => n30229, B1 => n26256, B2 => 
                           n30223, ZN => n28166);
   U21383 : AOI221_X1 port map( B1 => n30242, B2 => n22008, C1 => n30236, C2 =>
                           n9307, A => n28147, ZN => n28146);
   U21384 : OAI22_X1 port map( A1 => n26430, A2 => n30230, B1 => n26255, B2 => 
                           n30224, ZN => n28147);
   U21385 : AOI221_X1 port map( B1 => n30338, B2 => n21855, C1 => n30332, C2 =>
                           n9304, A => n28139, ZN => n28138);
   U21386 : OAI22_X1 port map( A1 => n8984, A2 => n30326, B1 => n9752, B2 => 
                           n30320, ZN => n28139);
   U21387 : AOI221_X1 port map( B1 => n30242, B2 => n22009, C1 => n30236, C2 =>
                           n9302, A => n28128, ZN => n28127);
   U21388 : OAI22_X1 port map( A1 => n26404, A2 => n30230, B1 => n26254, B2 => 
                           n30224, ZN => n28128);
   U21389 : AOI221_X1 port map( B1 => n30338, B2 => n21856, C1 => n30332, C2 =>
                           n9299, A => n28120, ZN => n28119);
   U21390 : OAI22_X1 port map( A1 => n8979, A2 => n30326, B1 => n9747, B2 => 
                           n30320, ZN => n28120);
   U21391 : AOI221_X1 port map( B1 => n30242, B2 => n22010, C1 => n30236, C2 =>
                           n9297, A => n28109, ZN => n28108);
   U21392 : OAI22_X1 port map( A1 => n26378, A2 => n30230, B1 => n26253, B2 => 
                           n30224, ZN => n28109);
   U21393 : AOI221_X1 port map( B1 => n30338, B2 => n21857, C1 => n30332, C2 =>
                           n9294, A => n28101, ZN => n28100);
   U21394 : OAI22_X1 port map( A1 => n8974, A2 => n30326, B1 => n9742, B2 => 
                           n30320, ZN => n28101);
   U21395 : AOI221_X1 port map( B1 => n30242, B2 => n22011, C1 => n30236, C2 =>
                           n9292, A => n28075, ZN => n28072);
   U21396 : OAI22_X1 port map( A1 => n26317, A2 => n30230, B1 => n26251, B2 => 
                           n30224, ZN => n28075);
   U21397 : AOI221_X1 port map( B1 => n30338, B2 => n21858, C1 => n30332, C2 =>
                           n9289, A => n28051, ZN => n28048);
   U21398 : OAI22_X1 port map( A1 => n8969, A2 => n30326, B1 => n9737, B2 => 
                           n30320, ZN => n28051);
   U21399 : AOI221_X1 port map( B1 => n30441, B2 => n21859, C1 => n30435, C2 =>
                           n9608, A => n28018, ZN => n28017);
   U21400 : OAI22_X1 port map( A1 => n26088, A2 => n30429, B1 => n26022, B2 => 
                           n30423, ZN => n28018);
   U21401 : AOI221_X1 port map( B1 => n30538, B2 => n21795, C1 => n30532, C2 =>
                           n9604, A => n27999, ZN => n27998);
   U21402 : OAI22_X1 port map( A1 => n9284, A2 => n30526, B1 => n25229, B2 => 
                           n30520, ZN => n27999);
   U21403 : AOI221_X1 port map( B1 => n30441, B2 => n21860, C1 => n30435, C2 =>
                           n9603, A => n27980, ZN => n27979);
   U21404 : OAI22_X1 port map( A1 => n26087, A2 => n30429, B1 => n26021, B2 => 
                           n30423, ZN => n27980);
   U21405 : AOI221_X1 port map( B1 => n30538, B2 => n21796, C1 => n30532, C2 =>
                           n9599, A => n27972, ZN => n27971);
   U21406 : OAI22_X1 port map( A1 => n9279, A2 => n30526, B1 => n25227, B2 => 
                           n30520, ZN => n27972);
   U21407 : AOI221_X1 port map( B1 => n30441, B2 => n21861, C1 => n30435, C2 =>
                           n9598, A => n27954, ZN => n27953);
   U21408 : OAI22_X1 port map( A1 => n26086, A2 => n30429, B1 => n26020, B2 => 
                           n30423, ZN => n27954);
   U21409 : AOI221_X1 port map( B1 => n30538, B2 => n21797, C1 => n30532, C2 =>
                           n9594, A => n27946, ZN => n27945);
   U21410 : OAI22_X1 port map( A1 => n9274, A2 => n30526, B1 => n25225, B2 => 
                           n30520, ZN => n27946);
   U21411 : AOI221_X1 port map( B1 => n30441, B2 => n21862, C1 => n30435, C2 =>
                           n9593, A => n27928, ZN => n27927);
   U21412 : OAI22_X1 port map( A1 => n26085, A2 => n30429, B1 => n26019, B2 => 
                           n30423, ZN => n27928);
   U21413 : AOI221_X1 port map( B1 => n30538, B2 => n21798, C1 => n30532, C2 =>
                           n9589, A => n27920, ZN => n27919);
   U21414 : OAI22_X1 port map( A1 => n9269, A2 => n30526, B1 => n25223, B2 => 
                           n30520, ZN => n27920);
   U21415 : AOI221_X1 port map( B1 => n30441, B2 => n21863, C1 => n30435, C2 =>
                           n9588, A => n27902, ZN => n27901);
   U21416 : OAI22_X1 port map( A1 => n26084, A2 => n30429, B1 => n26018, B2 => 
                           n30423, ZN => n27902);
   U21417 : AOI221_X1 port map( B1 => n30538, B2 => n21799, C1 => n30532, C2 =>
                           n9584, A => n27894, ZN => n27893);
   U21418 : OAI22_X1 port map( A1 => n9264, A2 => n30526, B1 => n25221, B2 => 
                           n30520, ZN => n27894);
   U21419 : AOI221_X1 port map( B1 => n30441, B2 => n21864, C1 => n30435, C2 =>
                           n9583, A => n27876, ZN => n27875);
   U21420 : OAI22_X1 port map( A1 => n26083, A2 => n30429, B1 => n26017, B2 => 
                           n30423, ZN => n27876);
   U21421 : AOI221_X1 port map( B1 => n30538, B2 => n21800, C1 => n30532, C2 =>
                           n9579, A => n27868, ZN => n27867);
   U21422 : OAI22_X1 port map( A1 => n9259, A2 => n30526, B1 => n25219, B2 => 
                           n30520, ZN => n27868);
   U21423 : AOI221_X1 port map( B1 => n30441, B2 => n21865, C1 => n30435, C2 =>
                           n9578, A => n27850, ZN => n27849);
   U21424 : OAI22_X1 port map( A1 => n26082, A2 => n30429, B1 => n26016, B2 => 
                           n30423, ZN => n27850);
   U21425 : AOI221_X1 port map( B1 => n30538, B2 => n21801, C1 => n30532, C2 =>
                           n9574, A => n27842, ZN => n27841);
   U21426 : OAI22_X1 port map( A1 => n9254, A2 => n30526, B1 => n25217, B2 => 
                           n30520, ZN => n27842);
   U21427 : AOI221_X1 port map( B1 => n30441, B2 => n21866, C1 => n30435, C2 =>
                           n9573, A => n27824, ZN => n27823);
   U21428 : OAI22_X1 port map( A1 => n26081, A2 => n30429, B1 => n26015, B2 => 
                           n30423, ZN => n27824);
   U21429 : AOI221_X1 port map( B1 => n30538, B2 => n21802, C1 => n30532, C2 =>
                           n9569, A => n27816, ZN => n27815);
   U21430 : OAI22_X1 port map( A1 => n9249, A2 => n30526, B1 => n25215, B2 => 
                           n30520, ZN => n27816);
   U21431 : AOI221_X1 port map( B1 => n30441, B2 => n21867, C1 => n30435, C2 =>
                           n9568, A => n27798, ZN => n27797);
   U21432 : OAI22_X1 port map( A1 => n26080, A2 => n30429, B1 => n26014, B2 => 
                           n30423, ZN => n27798);
   U21433 : AOI221_X1 port map( B1 => n30538, B2 => n21803, C1 => n30532, C2 =>
                           n9564, A => n27790, ZN => n27789);
   U21434 : OAI22_X1 port map( A1 => n9244, A2 => n30526, B1 => n25213, B2 => 
                           n30520, ZN => n27790);
   U21435 : AOI221_X1 port map( B1 => n30441, B2 => n21868, C1 => n30435, C2 =>
                           n9563, A => n27772, ZN => n27771);
   U21436 : OAI22_X1 port map( A1 => n26079, A2 => n30429, B1 => n26013, B2 => 
                           n30423, ZN => n27772);
   U21437 : AOI221_X1 port map( B1 => n30538, B2 => n21804, C1 => n30532, C2 =>
                           n9559, A => n27764, ZN => n27763);
   U21438 : OAI22_X1 port map( A1 => n9239, A2 => n30526, B1 => n25211, B2 => 
                           n30520, ZN => n27764);
   U21439 : AOI221_X1 port map( B1 => n30441, B2 => n21869, C1 => n30435, C2 =>
                           n9558, A => n27746, ZN => n27745);
   U21440 : OAI22_X1 port map( A1 => n26078, A2 => n30429, B1 => n26012, B2 => 
                           n30423, ZN => n27746);
   U21441 : AOI221_X1 port map( B1 => n30538, B2 => n21805, C1 => n30532, C2 =>
                           n9554, A => n27738, ZN => n27737);
   U21442 : OAI22_X1 port map( A1 => n9234, A2 => n30526, B1 => n25209, B2 => 
                           n30520, ZN => n27738);
   U21443 : AOI221_X1 port map( B1 => n30441, B2 => n21870, C1 => n30435, C2 =>
                           n9553, A => n27720, ZN => n27719);
   U21444 : OAI22_X1 port map( A1 => n26077, A2 => n30429, B1 => n26011, B2 => 
                           n30423, ZN => n27720);
   U21445 : AOI221_X1 port map( B1 => n30538, B2 => n21806, C1 => n30532, C2 =>
                           n9549, A => n27712, ZN => n27711);
   U21446 : OAI22_X1 port map( A1 => n9229, A2 => n30526, B1 => n9997, B2 => 
                           n30520, ZN => n27712);
   U21447 : AOI221_X1 port map( B1 => n30442, B2 => n21871, C1 => n30436, C2 =>
                           n9548, A => n27694, ZN => n27693);
   U21448 : OAI22_X1 port map( A1 => n26076, A2 => n30430, B1 => n26010, B2 => 
                           n30424, ZN => n27694);
   U21449 : AOI221_X1 port map( B1 => n30539, B2 => n21807, C1 => n30533, C2 =>
                           n9544, A => n27686, ZN => n27685);
   U21450 : OAI22_X1 port map( A1 => n9224, A2 => n30527, B1 => n9992, B2 => 
                           n30521, ZN => n27686);
   U21451 : AOI221_X1 port map( B1 => n30442, B2 => n21872, C1 => n30436, C2 =>
                           n9543, A => n27668, ZN => n27667);
   U21452 : OAI22_X1 port map( A1 => n26075, A2 => n30430, B1 => n26009, B2 => 
                           n30424, ZN => n27668);
   U21453 : AOI221_X1 port map( B1 => n30539, B2 => n21808, C1 => n30533, C2 =>
                           n9539, A => n27660, ZN => n27659);
   U21454 : OAI22_X1 port map( A1 => n9219, A2 => n30527, B1 => n9987, B2 => 
                           n30521, ZN => n27660);
   U21455 : AOI221_X1 port map( B1 => n30442, B2 => n21873, C1 => n30436, C2 =>
                           n9538, A => n27642, ZN => n27641);
   U21456 : OAI22_X1 port map( A1 => n26074, A2 => n30430, B1 => n26008, B2 => 
                           n30424, ZN => n27642);
   U21457 : AOI221_X1 port map( B1 => n30539, B2 => n21809, C1 => n30533, C2 =>
                           n9534, A => n27634, ZN => n27633);
   U21458 : OAI22_X1 port map( A1 => n9214, A2 => n30527, B1 => n9982, B2 => 
                           n30521, ZN => n27634);
   U21459 : AOI221_X1 port map( B1 => n30442, B2 => n21874, C1 => n30436, C2 =>
                           n9533, A => n27616, ZN => n27615);
   U21460 : OAI22_X1 port map( A1 => n26073, A2 => n30430, B1 => n26007, B2 => 
                           n30424, ZN => n27616);
   U21461 : AOI221_X1 port map( B1 => n30539, B2 => n21810, C1 => n30533, C2 =>
                           n9529, A => n27608, ZN => n27607);
   U21462 : OAI22_X1 port map( A1 => n9209, A2 => n30527, B1 => n9977, B2 => 
                           n30521, ZN => n27608);
   U21463 : AOI221_X1 port map( B1 => n30442, B2 => n21875, C1 => n30436, C2 =>
                           n9528, A => n27590, ZN => n27589);
   U21464 : OAI22_X1 port map( A1 => n26072, A2 => n30430, B1 => n26006, B2 => 
                           n30424, ZN => n27590);
   U21465 : AOI221_X1 port map( B1 => n30539, B2 => n21811, C1 => n30533, C2 =>
                           n9524, A => n27582, ZN => n27581);
   U21466 : OAI22_X1 port map( A1 => n9204, A2 => n30527, B1 => n9972, B2 => 
                           n30521, ZN => n27582);
   U21467 : AOI221_X1 port map( B1 => n30442, B2 => n21876, C1 => n30436, C2 =>
                           n9523, A => n27564, ZN => n27563);
   U21468 : OAI22_X1 port map( A1 => n26071, A2 => n30430, B1 => n26005, B2 => 
                           n30424, ZN => n27564);
   U21469 : AOI221_X1 port map( B1 => n30539, B2 => n21812, C1 => n30533, C2 =>
                           n9519, A => n27556, ZN => n27555);
   U21470 : OAI22_X1 port map( A1 => n9199, A2 => n30527, B1 => n9967, B2 => 
                           n30521, ZN => n27556);
   U21471 : AOI221_X1 port map( B1 => n30442, B2 => n21877, C1 => n30436, C2 =>
                           n9518, A => n27538, ZN => n27537);
   U21472 : OAI22_X1 port map( A1 => n26070, A2 => n30430, B1 => n26004, B2 => 
                           n30424, ZN => n27538);
   U21473 : AOI221_X1 port map( B1 => n30539, B2 => n21813, C1 => n30533, C2 =>
                           n9514, A => n27530, ZN => n27529);
   U21474 : OAI22_X1 port map( A1 => n9194, A2 => n30527, B1 => n9962, B2 => 
                           n30521, ZN => n27530);
   U21475 : AOI221_X1 port map( B1 => n30442, B2 => n21878, C1 => n30436, C2 =>
                           n9513, A => n27512, ZN => n27511);
   U21476 : OAI22_X1 port map( A1 => n26069, A2 => n30430, B1 => n26003, B2 => 
                           n30424, ZN => n27512);
   U21477 : AOI221_X1 port map( B1 => n30539, B2 => n21814, C1 => n30533, C2 =>
                           n9509, A => n27504, ZN => n27503);
   U21478 : OAI22_X1 port map( A1 => n9189, A2 => n30527, B1 => n9957, B2 => 
                           n30521, ZN => n27504);
   U21479 : AOI221_X1 port map( B1 => n30442, B2 => n21879, C1 => n30436, C2 =>
                           n9508, A => n27486, ZN => n27485);
   U21480 : OAI22_X1 port map( A1 => n26068, A2 => n30430, B1 => n26002, B2 => 
                           n30424, ZN => n27486);
   U21481 : AOI221_X1 port map( B1 => n30539, B2 => n21815, C1 => n30533, C2 =>
                           n9504, A => n27478, ZN => n27477);
   U21482 : OAI22_X1 port map( A1 => n9184, A2 => n30527, B1 => n9952, B2 => 
                           n30521, ZN => n27478);
   U21483 : AOI221_X1 port map( B1 => n30442, B2 => n21880, C1 => n30436, C2 =>
                           n9503, A => n27460, ZN => n27459);
   U21484 : OAI22_X1 port map( A1 => n26067, A2 => n30430, B1 => n26001, B2 => 
                           n30424, ZN => n27460);
   U21485 : AOI221_X1 port map( B1 => n30539, B2 => n21816, C1 => n30533, C2 =>
                           n9499, A => n27452, ZN => n27451);
   U21486 : OAI22_X1 port map( A1 => n9179, A2 => n30527, B1 => n9947, B2 => 
                           n30521, ZN => n27452);
   U21487 : AOI221_X1 port map( B1 => n30442, B2 => n21881, C1 => n30436, C2 =>
                           n9498, A => n27434, ZN => n27433);
   U21488 : OAI22_X1 port map( A1 => n26066, A2 => n30430, B1 => n26000, B2 => 
                           n30424, ZN => n27434);
   U21489 : AOI221_X1 port map( B1 => n30539, B2 => n21817, C1 => n30533, C2 =>
                           n9494, A => n27426, ZN => n27425);
   U21490 : OAI22_X1 port map( A1 => n9174, A2 => n30527, B1 => n9942, B2 => 
                           n30521, ZN => n27426);
   U21491 : AOI221_X1 port map( B1 => n30442, B2 => n21882, C1 => n30436, C2 =>
                           n9493, A => n27408, ZN => n27407);
   U21492 : OAI22_X1 port map( A1 => n26065, A2 => n30430, B1 => n25999, B2 => 
                           n30424, ZN => n27408);
   U21493 : AOI221_X1 port map( B1 => n30539, B2 => n21818, C1 => n30533, C2 =>
                           n9489, A => n27400, ZN => n27399);
   U21494 : OAI22_X1 port map( A1 => n9169, A2 => n30527, B1 => n9937, B2 => 
                           n30521, ZN => n27400);
   U21495 : AOI221_X1 port map( B1 => n30443, B2 => n21883, C1 => n30437, C2 =>
                           n9488, A => n27382, ZN => n27381);
   U21496 : OAI22_X1 port map( A1 => n26064, A2 => n30431, B1 => n25998, B2 => 
                           n30425, ZN => n27382);
   U21497 : AOI221_X1 port map( B1 => n30540, B2 => n21819, C1 => n30534, C2 =>
                           n9484, A => n27374, ZN => n27373);
   U21498 : OAI22_X1 port map( A1 => n9164, A2 => n30528, B1 => n9932, B2 => 
                           n30522, ZN => n27374);
   U21499 : AOI221_X1 port map( B1 => n30540, B2 => n21820, C1 => n30534, C2 =>
                           n9479, A => n27348, ZN => n27347);
   U21500 : OAI22_X1 port map( A1 => n9159, A2 => n30528, B1 => n9927, B2 => 
                           n30522, ZN => n27348);
   U21501 : AOI221_X1 port map( B1 => n30443, B2 => n21884, C1 => n30437, C2 =>
                           n9483, A => n27356, ZN => n27355);
   U21502 : OAI22_X1 port map( A1 => n26063, A2 => n30431, B1 => n25997, B2 => 
                           n30425, ZN => n27356);
   U21503 : AOI221_X1 port map( B1 => n30540, B2 => n21821, C1 => n30534, C2 =>
                           n9474, A => n27322, ZN => n27321);
   U21504 : OAI22_X1 port map( A1 => n9154, A2 => n30528, B1 => n9922, B2 => 
                           n30522, ZN => n27322);
   U21505 : AOI221_X1 port map( B1 => n30443, B2 => n21885, C1 => n30437, C2 =>
                           n9478, A => n27330, ZN => n27329);
   U21506 : OAI22_X1 port map( A1 => n26062, A2 => n30431, B1 => n25996, B2 => 
                           n30425, ZN => n27330);
   U21507 : AOI221_X1 port map( B1 => n30540, B2 => n21822, C1 => n30534, C2 =>
                           n9469, A => n27296, ZN => n27295);
   U21508 : OAI22_X1 port map( A1 => n9149, A2 => n30528, B1 => n9917, B2 => 
                           n30522, ZN => n27296);
   U21509 : AOI221_X1 port map( B1 => n30443, B2 => n21886, C1 => n30437, C2 =>
                           n9473, A => n27304, ZN => n27303);
   U21510 : OAI22_X1 port map( A1 => n26061, A2 => n30431, B1 => n25995, B2 => 
                           n30425, ZN => n27304);
   U21511 : AOI221_X1 port map( B1 => n30540, B2 => n21823, C1 => n30534, C2 =>
                           n9464, A => n27270, ZN => n27269);
   U21512 : OAI22_X1 port map( A1 => n9144, A2 => n30528, B1 => n9912, B2 => 
                           n30522, ZN => n27270);
   U21513 : AOI221_X1 port map( B1 => n30443, B2 => n21887, C1 => n30437, C2 =>
                           n9468, A => n27278, ZN => n27277);
   U21514 : OAI22_X1 port map( A1 => n26060, A2 => n30431, B1 => n25994, B2 => 
                           n30425, ZN => n27278);
   U21515 : AOI221_X1 port map( B1 => n30540, B2 => n21824, C1 => n30534, C2 =>
                           n9459, A => n27244, ZN => n27243);
   U21516 : OAI22_X1 port map( A1 => n9139, A2 => n30528, B1 => n9907, B2 => 
                           n30522, ZN => n27244);
   U21517 : AOI221_X1 port map( B1 => n30443, B2 => n21888, C1 => n30437, C2 =>
                           n9463, A => n27252, ZN => n27251);
   U21518 : OAI22_X1 port map( A1 => n26059, A2 => n30431, B1 => n25993, B2 => 
                           n30425, ZN => n27252);
   U21519 : AOI221_X1 port map( B1 => n30540, B2 => n21825, C1 => n30534, C2 =>
                           n9454, A => n27218, ZN => n27217);
   U21520 : OAI22_X1 port map( A1 => n9134, A2 => n30528, B1 => n9902, B2 => 
                           n30522, ZN => n27218);
   U21521 : AOI221_X1 port map( B1 => n30443, B2 => n21889, C1 => n30437, C2 =>
                           n9458, A => n27226, ZN => n27225);
   U21522 : OAI22_X1 port map( A1 => n26058, A2 => n30431, B1 => n25992, B2 => 
                           n30425, ZN => n27226);
   U21523 : AOI221_X1 port map( B1 => n30540, B2 => n21826, C1 => n30534, C2 =>
                           n9449, A => n27192, ZN => n27191);
   U21524 : OAI22_X1 port map( A1 => n9129, A2 => n30528, B1 => n9897, B2 => 
                           n30522, ZN => n27192);
   U21525 : AOI221_X1 port map( B1 => n30443, B2 => n21890, C1 => n30437, C2 =>
                           n9453, A => n27200, ZN => n27199);
   U21526 : OAI22_X1 port map( A1 => n26057, A2 => n30431, B1 => n25991, B2 => 
                           n30425, ZN => n27200);
   U21527 : AOI221_X1 port map( B1 => n30540, B2 => n21827, C1 => n30534, C2 =>
                           n9444, A => n27166, ZN => n27165);
   U21528 : OAI22_X1 port map( A1 => n9124, A2 => n30528, B1 => n9892, B2 => 
                           n30522, ZN => n27166);
   U21529 : AOI221_X1 port map( B1 => n30443, B2 => n21891, C1 => n30437, C2 =>
                           n9448, A => n27174, ZN => n27173);
   U21530 : OAI22_X1 port map( A1 => n26056, A2 => n30431, B1 => n25990, B2 => 
                           n30425, ZN => n27174);
   U21531 : AOI221_X1 port map( B1 => n30540, B2 => n21828, C1 => n30534, C2 =>
                           n9439, A => n27140, ZN => n27139);
   U21532 : OAI22_X1 port map( A1 => n9119, A2 => n30528, B1 => n9887, B2 => 
                           n30522, ZN => n27140);
   U21533 : AOI221_X1 port map( B1 => n30443, B2 => n21892, C1 => n30437, C2 =>
                           n9443, A => n27148, ZN => n27147);
   U21534 : OAI22_X1 port map( A1 => n26055, A2 => n30431, B1 => n25989, B2 => 
                           n30425, ZN => n27148);
   U21535 : AOI221_X1 port map( B1 => n30540, B2 => n21829, C1 => n30534, C2 =>
                           n9434, A => n27114, ZN => n27113);
   U21536 : OAI22_X1 port map( A1 => n9114, A2 => n30528, B1 => n9882, B2 => 
                           n30522, ZN => n27114);
   U21537 : AOI221_X1 port map( B1 => n30443, B2 => n21893, C1 => n30437, C2 =>
                           n9438, A => n27122, ZN => n27121);
   U21538 : OAI22_X1 port map( A1 => n26054, A2 => n30431, B1 => n25988, B2 => 
                           n30425, ZN => n27122);
   U21539 : AOI221_X1 port map( B1 => n30540, B2 => n21830, C1 => n30534, C2 =>
                           n9429, A => n27088, ZN => n27087);
   U21540 : OAI22_X1 port map( A1 => n9109, A2 => n30528, B1 => n9877, B2 => 
                           n30522, ZN => n27088);
   U21541 : AOI221_X1 port map( B1 => n30443, B2 => n21894, C1 => n30437, C2 =>
                           n9433, A => n27096, ZN => n27095);
   U21542 : OAI22_X1 port map( A1 => n26053, A2 => n30431, B1 => n25987, B2 => 
                           n30425, ZN => n27096);
   U21543 : AOI221_X1 port map( B1 => n30541, B2 => n21831, C1 => n30535, C2 =>
                           n9424, A => n27062, ZN => n27061);
   U21544 : OAI22_X1 port map( A1 => n9104, A2 => n30529, B1 => n9872, B2 => 
                           n30523, ZN => n27062);
   U21545 : AOI221_X1 port map( B1 => n30444, B2 => n21895, C1 => n30438, C2 =>
                           n9428, A => n27070, ZN => n27069);
   U21546 : OAI22_X1 port map( A1 => n26052, A2 => n30432, B1 => n25986, B2 => 
                           n30426, ZN => n27070);
   U21547 : AOI221_X1 port map( B1 => n30541, B2 => n21832, C1 => n30535, C2 =>
                           n9419, A => n27036, ZN => n27035);
   U21548 : OAI22_X1 port map( A1 => n9099, A2 => n30529, B1 => n9867, B2 => 
                           n30523, ZN => n27036);
   U21549 : AOI221_X1 port map( B1 => n30444, B2 => n21896, C1 => n30438, C2 =>
                           n9423, A => n27044, ZN => n27043);
   U21550 : OAI22_X1 port map( A1 => n26051, A2 => n30432, B1 => n25985, B2 => 
                           n30426, ZN => n27044);
   U21551 : AOI221_X1 port map( B1 => n30541, B2 => n21833, C1 => n30535, C2 =>
                           n9414, A => n27010, ZN => n27009);
   U21552 : OAI22_X1 port map( A1 => n9094, A2 => n30529, B1 => n9862, B2 => 
                           n30523, ZN => n27010);
   U21553 : AOI221_X1 port map( B1 => n30444, B2 => n21897, C1 => n30438, C2 =>
                           n9418, A => n27018, ZN => n27017);
   U21554 : OAI22_X1 port map( A1 => n26050, A2 => n30432, B1 => n25984, B2 => 
                           n30426, ZN => n27018);
   U21555 : AOI221_X1 port map( B1 => n30541, B2 => n21834, C1 => n30535, C2 =>
                           n9409, A => n26984, ZN => n26983);
   U21556 : OAI22_X1 port map( A1 => n9089, A2 => n30529, B1 => n9857, B2 => 
                           n30523, ZN => n26984);
   U21557 : AOI221_X1 port map( B1 => n30444, B2 => n21898, C1 => n30438, C2 =>
                           n9413, A => n26992, ZN => n26991);
   U21558 : OAI22_X1 port map( A1 => n26049, A2 => n30432, B1 => n25983, B2 => 
                           n30426, ZN => n26992);
   U21559 : AOI221_X1 port map( B1 => n30541, B2 => n21835, C1 => n30535, C2 =>
                           n9404, A => n26958, ZN => n26957);
   U21560 : OAI22_X1 port map( A1 => n9084, A2 => n30529, B1 => n9852, B2 => 
                           n30523, ZN => n26958);
   U21561 : AOI221_X1 port map( B1 => n30444, B2 => n21899, C1 => n30438, C2 =>
                           n9408, A => n26966, ZN => n26965);
   U21562 : OAI22_X1 port map( A1 => n26048, A2 => n30432, B1 => n25982, B2 => 
                           n30426, ZN => n26966);
   U21563 : AOI221_X1 port map( B1 => n30541, B2 => n21836, C1 => n30535, C2 =>
                           n9399, A => n26932, ZN => n26931);
   U21564 : OAI22_X1 port map( A1 => n9079, A2 => n30529, B1 => n9847, B2 => 
                           n30523, ZN => n26932);
   U21565 : AOI221_X1 port map( B1 => n30444, B2 => n21900, C1 => n30438, C2 =>
                           n9403, A => n26940, ZN => n26939);
   U21566 : OAI22_X1 port map( A1 => n26047, A2 => n30432, B1 => n25981, B2 => 
                           n30426, ZN => n26940);
   U21567 : AOI221_X1 port map( B1 => n30541, B2 => n21837, C1 => n30535, C2 =>
                           n9394, A => n26906, ZN => n26905);
   U21568 : OAI22_X1 port map( A1 => n9074, A2 => n30529, B1 => n9842, B2 => 
                           n30523, ZN => n26906);
   U21569 : AOI221_X1 port map( B1 => n30444, B2 => n21901, C1 => n30438, C2 =>
                           n9398, A => n26914, ZN => n26913);
   U21570 : OAI22_X1 port map( A1 => n26046, A2 => n30432, B1 => n25980, B2 => 
                           n30426, ZN => n26914);
   U21571 : AOI221_X1 port map( B1 => n30541, B2 => n21838, C1 => n30535, C2 =>
                           n9389, A => n26880, ZN => n26879);
   U21572 : OAI22_X1 port map( A1 => n9069, A2 => n30529, B1 => n9837, B2 => 
                           n30523, ZN => n26880);
   U21573 : AOI221_X1 port map( B1 => n30444, B2 => n21902, C1 => n30438, C2 =>
                           n9393, A => n26888, ZN => n26887);
   U21574 : OAI22_X1 port map( A1 => n26045, A2 => n30432, B1 => n25979, B2 => 
                           n30426, ZN => n26888);
   U21575 : AOI221_X1 port map( B1 => n30541, B2 => n21839, C1 => n30535, C2 =>
                           n9384, A => n26854, ZN => n26853);
   U21576 : OAI22_X1 port map( A1 => n9064, A2 => n30529, B1 => n9832, B2 => 
                           n30523, ZN => n26854);
   U21577 : AOI221_X1 port map( B1 => n30444, B2 => n21903, C1 => n30438, C2 =>
                           n9388, A => n26862, ZN => n26861);
   U21578 : OAI22_X1 port map( A1 => n26044, A2 => n30432, B1 => n25978, B2 => 
                           n30426, ZN => n26862);
   U21579 : AOI221_X1 port map( B1 => n30541, B2 => n21840, C1 => n30535, C2 =>
                           n9379, A => n26828, ZN => n26827);
   U21580 : OAI22_X1 port map( A1 => n9059, A2 => n30529, B1 => n9827, B2 => 
                           n30523, ZN => n26828);
   U21581 : AOI221_X1 port map( B1 => n30444, B2 => n21904, C1 => n30438, C2 =>
                           n9383, A => n26836, ZN => n26835);
   U21582 : OAI22_X1 port map( A1 => n26043, A2 => n30432, B1 => n25977, B2 => 
                           n30426, ZN => n26836);
   U21583 : AOI221_X1 port map( B1 => n30541, B2 => n21841, C1 => n30535, C2 =>
                           n9374, A => n26802, ZN => n26801);
   U21584 : OAI22_X1 port map( A1 => n9054, A2 => n30529, B1 => n9822, B2 => 
                           n30523, ZN => n26802);
   U21585 : AOI221_X1 port map( B1 => n30444, B2 => n21905, C1 => n30438, C2 =>
                           n9378, A => n26810, ZN => n26809);
   U21586 : OAI22_X1 port map( A1 => n26042, A2 => n30432, B1 => n25976, B2 => 
                           n30426, ZN => n26810);
   U21587 : AOI221_X1 port map( B1 => n30541, B2 => n21842, C1 => n30535, C2 =>
                           n9369, A => n26776, ZN => n26775);
   U21588 : OAI22_X1 port map( A1 => n9049, A2 => n30529, B1 => n9817, B2 => 
                           n30523, ZN => n26776);
   U21589 : AOI221_X1 port map( B1 => n30444, B2 => n21906, C1 => n30438, C2 =>
                           n9373, A => n26784, ZN => n26783);
   U21590 : OAI22_X1 port map( A1 => n26041, A2 => n30432, B1 => n25975, B2 => 
                           n30426, ZN => n26784);
   U21591 : AOI221_X1 port map( B1 => n30542, B2 => n21843, C1 => n30536, C2 =>
                           n9364, A => n26750, ZN => n26749);
   U21592 : OAI22_X1 port map( A1 => n9044, A2 => n30530, B1 => n9812, B2 => 
                           n30524, ZN => n26750);
   U21593 : AOI221_X1 port map( B1 => n30445, B2 => n21907, C1 => n30439, C2 =>
                           n9368, A => n26758, ZN => n26757);
   U21594 : OAI22_X1 port map( A1 => n26040, A2 => n30433, B1 => n25974, B2 => 
                           n30427, ZN => n26758);
   U21595 : AOI221_X1 port map( B1 => n30542, B2 => n21844, C1 => n30536, C2 =>
                           n9359, A => n26724, ZN => n26723);
   U21596 : OAI22_X1 port map( A1 => n9039, A2 => n30530, B1 => n9807, B2 => 
                           n30524, ZN => n26724);
   U21597 : AOI221_X1 port map( B1 => n30445, B2 => n21908, C1 => n30439, C2 =>
                           n9363, A => n26732, ZN => n26731);
   U21598 : OAI22_X1 port map( A1 => n26039, A2 => n30433, B1 => n25973, B2 => 
                           n30427, ZN => n26732);
   U21599 : AOI221_X1 port map( B1 => n30542, B2 => n21845, C1 => n30536, C2 =>
                           n9354, A => n26698, ZN => n26697);
   U21600 : OAI22_X1 port map( A1 => n9034, A2 => n30530, B1 => n9802, B2 => 
                           n30524, ZN => n26698);
   U21601 : AOI221_X1 port map( B1 => n30445, B2 => n21909, C1 => n30439, C2 =>
                           n9358, A => n26706, ZN => n26705);
   U21602 : OAI22_X1 port map( A1 => n26038, A2 => n30433, B1 => n25972, B2 => 
                           n30427, ZN => n26706);
   U21603 : AOI221_X1 port map( B1 => n30542, B2 => n21846, C1 => n30536, C2 =>
                           n9349, A => n26672, ZN => n26671);
   U21604 : OAI22_X1 port map( A1 => n9029, A2 => n30530, B1 => n9797, B2 => 
                           n30524, ZN => n26672);
   U21605 : AOI221_X1 port map( B1 => n30445, B2 => n21910, C1 => n30439, C2 =>
                           n9353, A => n26680, ZN => n26679);
   U21606 : OAI22_X1 port map( A1 => n26037, A2 => n30433, B1 => n25971, B2 => 
                           n30427, ZN => n26680);
   U21607 : AOI221_X1 port map( B1 => n30542, B2 => n21847, C1 => n30536, C2 =>
                           n9344, A => n26646, ZN => n26645);
   U21608 : OAI22_X1 port map( A1 => n9024, A2 => n30530, B1 => n9792, B2 => 
                           n30524, ZN => n26646);
   U21609 : AOI221_X1 port map( B1 => n30445, B2 => n21911, C1 => n30439, C2 =>
                           n9348, A => n26654, ZN => n26653);
   U21610 : OAI22_X1 port map( A1 => n26036, A2 => n30433, B1 => n25970, B2 => 
                           n30427, ZN => n26654);
   U21611 : AOI221_X1 port map( B1 => n30542, B2 => n21848, C1 => n30536, C2 =>
                           n9339, A => n26620, ZN => n26619);
   U21612 : OAI22_X1 port map( A1 => n9019, A2 => n30530, B1 => n9787, B2 => 
                           n30524, ZN => n26620);
   U21613 : AOI221_X1 port map( B1 => n30445, B2 => n21912, C1 => n30439, C2 =>
                           n9343, A => n26628, ZN => n26627);
   U21614 : OAI22_X1 port map( A1 => n26035, A2 => n30433, B1 => n25969, B2 => 
                           n30427, ZN => n26628);
   U21615 : AOI221_X1 port map( B1 => n30542, B2 => n21849, C1 => n30536, C2 =>
                           n9334, A => n26594, ZN => n26593);
   U21616 : OAI22_X1 port map( A1 => n9014, A2 => n30530, B1 => n9782, B2 => 
                           n30524, ZN => n26594);
   U21617 : AOI221_X1 port map( B1 => n30445, B2 => n21913, C1 => n30439, C2 =>
                           n9338, A => n26602, ZN => n26601);
   U21618 : OAI22_X1 port map( A1 => n26034, A2 => n30433, B1 => n25968, B2 => 
                           n30427, ZN => n26602);
   U21619 : AOI221_X1 port map( B1 => n30542, B2 => n21850, C1 => n30536, C2 =>
                           n9329, A => n26568, ZN => n26567);
   U21620 : OAI22_X1 port map( A1 => n9009, A2 => n30530, B1 => n9777, B2 => 
                           n30524, ZN => n26568);
   U21621 : AOI221_X1 port map( B1 => n30445, B2 => n21914, C1 => n30439, C2 =>
                           n9333, A => n26576, ZN => n26575);
   U21622 : OAI22_X1 port map( A1 => n26033, A2 => n30433, B1 => n25967, B2 => 
                           n30427, ZN => n26576);
   U21623 : AOI221_X1 port map( B1 => n30542, B2 => n21851, C1 => n30536, C2 =>
                           n9324, A => n26542, ZN => n26541);
   U21624 : OAI22_X1 port map( A1 => n9004, A2 => n30530, B1 => n9772, B2 => 
                           n30524, ZN => n26542);
   U21625 : AOI221_X1 port map( B1 => n30445, B2 => n21915, C1 => n30439, C2 =>
                           n9328, A => n26550, ZN => n26549);
   U21626 : OAI22_X1 port map( A1 => n26032, A2 => n30433, B1 => n25966, B2 => 
                           n30427, ZN => n26550);
   U21627 : AOI221_X1 port map( B1 => n30542, B2 => n21852, C1 => n30536, C2 =>
                           n9319, A => n26516, ZN => n26515);
   U21628 : OAI22_X1 port map( A1 => n8999, A2 => n30530, B1 => n9767, B2 => 
                           n30524, ZN => n26516);
   U21629 : AOI221_X1 port map( B1 => n30445, B2 => n21916, C1 => n30439, C2 =>
                           n9323, A => n26524, ZN => n26523);
   U21630 : OAI22_X1 port map( A1 => n26031, A2 => n30433, B1 => n25965, B2 => 
                           n30427, ZN => n26524);
   U21631 : AOI221_X1 port map( B1 => n30542, B2 => n21853, C1 => n30536, C2 =>
                           n9314, A => n26490, ZN => n26489);
   U21632 : OAI22_X1 port map( A1 => n8994, A2 => n30530, B1 => n9762, B2 => 
                           n30524, ZN => n26490);
   U21633 : AOI221_X1 port map( B1 => n30445, B2 => n21917, C1 => n30439, C2 =>
                           n9318, A => n26498, ZN => n26497);
   U21634 : OAI22_X1 port map( A1 => n26030, A2 => n30433, B1 => n25964, B2 => 
                           n30427, ZN => n26498);
   U21635 : AOI221_X1 port map( B1 => n30542, B2 => n21854, C1 => n30536, C2 =>
                           n9309, A => n26464, ZN => n26463);
   U21636 : OAI22_X1 port map( A1 => n8989, A2 => n30530, B1 => n9757, B2 => 
                           n30524, ZN => n26464);
   U21637 : AOI221_X1 port map( B1 => n30445, B2 => n21918, C1 => n30439, C2 =>
                           n9313, A => n26472, ZN => n26471);
   U21638 : OAI22_X1 port map( A1 => n26029, A2 => n30433, B1 => n25963, B2 => 
                           n30427, ZN => n26472);
   U21639 : AOI221_X1 port map( B1 => n30543, B2 => n21855, C1 => n30537, C2 =>
                           n9304, A => n26438, ZN => n26437);
   U21640 : OAI22_X1 port map( A1 => n8984, A2 => n30531, B1 => n9752, B2 => 
                           n30525, ZN => n26438);
   U21641 : AOI221_X1 port map( B1 => n30543, B2 => n21856, C1 => n30537, C2 =>
                           n9299, A => n26412, ZN => n26411);
   U21642 : OAI22_X1 port map( A1 => n8979, A2 => n30531, B1 => n9747, B2 => 
                           n30525, ZN => n26412);
   U21643 : AOI221_X1 port map( B1 => n30543, B2 => n21857, C1 => n30537, C2 =>
                           n9294, A => n26386, ZN => n26385);
   U21644 : OAI22_X1 port map( A1 => n8974, A2 => n30531, B1 => n9742, B2 => 
                           n30525, ZN => n26386);
   U21645 : AOI221_X1 port map( B1 => n30543, B2 => n21858, C1 => n30537, C2 =>
                           n9289, A => n26330, ZN => n26327);
   U21646 : OAI22_X1 port map( A1 => n8969, A2 => n30531, B1 => n9737, B2 => 
                           n30525, ZN => n26330);
   U21647 : NOR3_X1 port map( A1 => n25152, A2 => ADD_WR(4), A3 => n25806, ZN 
                           => n25454);
   U21648 : AOI221_X1 port map( B1 => n30309, B2 => n22065, C1 => n30303, C2 =>
                           n9605, A => n29285, ZN => n29278);
   U21649 : OAI22_X1 port map( A1 => n9285, A2 => n30297, B1 => n25381, B2 => 
                           n30291, ZN => n29285);
   U21650 : AOI221_X1 port map( B1 => n30309, B2 => n22066, C1 => n30303, C2 =>
                           n9600, A => n29261, ZN => n29258);
   U21651 : OAI22_X1 port map( A1 => n9280, A2 => n30297, B1 => n25380, B2 => 
                           n30291, ZN => n29261);
   U21652 : AOI221_X1 port map( B1 => n30309, B2 => n22067, C1 => n30303, C2 =>
                           n9595, A => n29242, ZN => n29239);
   U21653 : OAI22_X1 port map( A1 => n9275, A2 => n30297, B1 => n25379, B2 => 
                           n30291, ZN => n29242);
   U21654 : AOI221_X1 port map( B1 => n30309, B2 => n22068, C1 => n30303, C2 =>
                           n9590, A => n29223, ZN => n29220);
   U21655 : OAI22_X1 port map( A1 => n9270, A2 => n30297, B1 => n25378, B2 => 
                           n30291, ZN => n29223);
   U21656 : AOI221_X1 port map( B1 => n30309, B2 => n22069, C1 => n30303, C2 =>
                           n9585, A => n29204, ZN => n29201);
   U21657 : OAI22_X1 port map( A1 => n9265, A2 => n30297, B1 => n25377, B2 => 
                           n30291, ZN => n29204);
   U21658 : AOI221_X1 port map( B1 => n30309, B2 => n22070, C1 => n30303, C2 =>
                           n9580, A => n29185, ZN => n29182);
   U21659 : OAI22_X1 port map( A1 => n9260, A2 => n30297, B1 => n25376, B2 => 
                           n30291, ZN => n29185);
   U21660 : AOI221_X1 port map( B1 => n30309, B2 => n22071, C1 => n30303, C2 =>
                           n9575, A => n29166, ZN => n29163);
   U21661 : OAI22_X1 port map( A1 => n9255, A2 => n30297, B1 => n25375, B2 => 
                           n30291, ZN => n29166);
   U21662 : AOI221_X1 port map( B1 => n30309, B2 => n22072, C1 => n30303, C2 =>
                           n9570, A => n29147, ZN => n29144);
   U21663 : OAI22_X1 port map( A1 => n9250, A2 => n30297, B1 => n25374, B2 => 
                           n30291, ZN => n29147);
   U21664 : AOI221_X1 port map( B1 => n30309, B2 => n22073, C1 => n30303, C2 =>
                           n9565, A => n29128, ZN => n29125);
   U21665 : OAI22_X1 port map( A1 => n9245, A2 => n30297, B1 => n25373, B2 => 
                           n30291, ZN => n29128);
   U21666 : AOI221_X1 port map( B1 => n30309, B2 => n22074, C1 => n30303, C2 =>
                           n9560, A => n29109, ZN => n29106);
   U21667 : OAI22_X1 port map( A1 => n9240, A2 => n30297, B1 => n25372, B2 => 
                           n30291, ZN => n29109);
   U21668 : AOI221_X1 port map( B1 => n30309, B2 => n22075, C1 => n30303, C2 =>
                           n9555, A => n29090, ZN => n29087);
   U21669 : OAI22_X1 port map( A1 => n9235, A2 => n30297, B1 => n25371, B2 => 
                           n30291, ZN => n29090);
   U21670 : AOI221_X1 port map( B1 => n30309, B2 => n22016, C1 => n30303, C2 =>
                           n9550, A => n29071, ZN => n29068);
   U21671 : OAI22_X1 port map( A1 => n9230, A2 => n30297, B1 => n9998, B2 => 
                           n30291, ZN => n29071);
   U21672 : AOI221_X1 port map( B1 => n30310, B2 => n22017, C1 => n30304, C2 =>
                           n9545, A => n29052, ZN => n29049);
   U21673 : OAI22_X1 port map( A1 => n9225, A2 => n30298, B1 => n9993, B2 => 
                           n30292, ZN => n29052);
   U21674 : AOI221_X1 port map( B1 => n30310, B2 => n22018, C1 => n30304, C2 =>
                           n9540, A => n29033, ZN => n29030);
   U21675 : OAI22_X1 port map( A1 => n9220, A2 => n30298, B1 => n9988, B2 => 
                           n30292, ZN => n29033);
   U21676 : AOI221_X1 port map( B1 => n30310, B2 => n22019, C1 => n30304, C2 =>
                           n9535, A => n29014, ZN => n29011);
   U21677 : OAI22_X1 port map( A1 => n9215, A2 => n30298, B1 => n9983, B2 => 
                           n30292, ZN => n29014);
   U21678 : AOI221_X1 port map( B1 => n30310, B2 => n22020, C1 => n30304, C2 =>
                           n9530, A => n28995, ZN => n28992);
   U21679 : OAI22_X1 port map( A1 => n9210, A2 => n30298, B1 => n9978, B2 => 
                           n30292, ZN => n28995);
   U21680 : AOI221_X1 port map( B1 => n30310, B2 => n22021, C1 => n30304, C2 =>
                           n9525, A => n28976, ZN => n28973);
   U21681 : OAI22_X1 port map( A1 => n9205, A2 => n30298, B1 => n9973, B2 => 
                           n30292, ZN => n28976);
   U21682 : AOI221_X1 port map( B1 => n30310, B2 => n22022, C1 => n30304, C2 =>
                           n9520, A => n28957, ZN => n28954);
   U21683 : OAI22_X1 port map( A1 => n9200, A2 => n30298, B1 => n9968, B2 => 
                           n30292, ZN => n28957);
   U21684 : AOI221_X1 port map( B1 => n30310, B2 => n22023, C1 => n30304, C2 =>
                           n9515, A => n28938, ZN => n28935);
   U21685 : OAI22_X1 port map( A1 => n9195, A2 => n30298, B1 => n9963, B2 => 
                           n30292, ZN => n28938);
   U21686 : AOI221_X1 port map( B1 => n30310, B2 => n22024, C1 => n30304, C2 =>
                           n9510, A => n28919, ZN => n28916);
   U21687 : OAI22_X1 port map( A1 => n9190, A2 => n30298, B1 => n9958, B2 => 
                           n30292, ZN => n28919);
   U21688 : AOI221_X1 port map( B1 => n30310, B2 => n22025, C1 => n30304, C2 =>
                           n9505, A => n28900, ZN => n28897);
   U21689 : OAI22_X1 port map( A1 => n9185, A2 => n30298, B1 => n9953, B2 => 
                           n30292, ZN => n28900);
   U21690 : AOI221_X1 port map( B1 => n30310, B2 => n22026, C1 => n30304, C2 =>
                           n9500, A => n28881, ZN => n28878);
   U21691 : OAI22_X1 port map( A1 => n9180, A2 => n30298, B1 => n9948, B2 => 
                           n30292, ZN => n28881);
   U21692 : AOI221_X1 port map( B1 => n30310, B2 => n22027, C1 => n30304, C2 =>
                           n9495, A => n28862, ZN => n28859);
   U21693 : OAI22_X1 port map( A1 => n9175, A2 => n30298, B1 => n9943, B2 => 
                           n30292, ZN => n28862);
   U21694 : AOI221_X1 port map( B1 => n30310, B2 => n22028, C1 => n30304, C2 =>
                           n9490, A => n28843, ZN => n28840);
   U21695 : OAI22_X1 port map( A1 => n9170, A2 => n30298, B1 => n9938, B2 => 
                           n30292, ZN => n28843);
   U21696 : AOI221_X1 port map( B1 => n30311, B2 => n22029, C1 => n30305, C2 =>
                           n9485, A => n28824, ZN => n28821);
   U21697 : OAI22_X1 port map( A1 => n9165, A2 => n30299, B1 => n9933, B2 => 
                           n30293, ZN => n28824);
   U21698 : AOI221_X1 port map( B1 => n30311, B2 => n22030, C1 => n30305, C2 =>
                           n9480, A => n28805, ZN => n28802);
   U21699 : OAI22_X1 port map( A1 => n9160, A2 => n30299, B1 => n9928, B2 => 
                           n30293, ZN => n28805);
   U21700 : AOI221_X1 port map( B1 => n30311, B2 => n22031, C1 => n30305, C2 =>
                           n9475, A => n28786, ZN => n28783);
   U21701 : OAI22_X1 port map( A1 => n9155, A2 => n30299, B1 => n9923, B2 => 
                           n30293, ZN => n28786);
   U21702 : AOI221_X1 port map( B1 => n30311, B2 => n22032, C1 => n30305, C2 =>
                           n9470, A => n28767, ZN => n28764);
   U21703 : OAI22_X1 port map( A1 => n9150, A2 => n30299, B1 => n9918, B2 => 
                           n30293, ZN => n28767);
   U21704 : AOI221_X1 port map( B1 => n30311, B2 => n22033, C1 => n30305, C2 =>
                           n9465, A => n28748, ZN => n28745);
   U21705 : OAI22_X1 port map( A1 => n9145, A2 => n30299, B1 => n9913, B2 => 
                           n30293, ZN => n28748);
   U21706 : AOI221_X1 port map( B1 => n30311, B2 => n22034, C1 => n30305, C2 =>
                           n9460, A => n28729, ZN => n28726);
   U21707 : OAI22_X1 port map( A1 => n9140, A2 => n30299, B1 => n9908, B2 => 
                           n30293, ZN => n28729);
   U21708 : AOI221_X1 port map( B1 => n30311, B2 => n22035, C1 => n30305, C2 =>
                           n9455, A => n28710, ZN => n28707);
   U21709 : OAI22_X1 port map( A1 => n9135, A2 => n30299, B1 => n9903, B2 => 
                           n30293, ZN => n28710);
   U21710 : AOI221_X1 port map( B1 => n30311, B2 => n22036, C1 => n30305, C2 =>
                           n9450, A => n28691, ZN => n28688);
   U21711 : OAI22_X1 port map( A1 => n9130, A2 => n30299, B1 => n9898, B2 => 
                           n30293, ZN => n28691);
   U21712 : AOI221_X1 port map( B1 => n30311, B2 => n22037, C1 => n30305, C2 =>
                           n9445, A => n28672, ZN => n28669);
   U21713 : OAI22_X1 port map( A1 => n9125, A2 => n30299, B1 => n9893, B2 => 
                           n30293, ZN => n28672);
   U21714 : AOI221_X1 port map( B1 => n30311, B2 => n22038, C1 => n30305, C2 =>
                           n9440, A => n28653, ZN => n28650);
   U21715 : OAI22_X1 port map( A1 => n9120, A2 => n30299, B1 => n9888, B2 => 
                           n30293, ZN => n28653);
   U21716 : AOI221_X1 port map( B1 => n30311, B2 => n22039, C1 => n30305, C2 =>
                           n9435, A => n28634, ZN => n28631);
   U21717 : OAI22_X1 port map( A1 => n9115, A2 => n30299, B1 => n9883, B2 => 
                           n30293, ZN => n28634);
   U21718 : AOI221_X1 port map( B1 => n30311, B2 => n22040, C1 => n30305, C2 =>
                           n9430, A => n28615, ZN => n28612);
   U21719 : OAI22_X1 port map( A1 => n9110, A2 => n30299, B1 => n9878, B2 => 
                           n30293, ZN => n28615);
   U21720 : AOI221_X1 port map( B1 => n30312, B2 => n22041, C1 => n30306, C2 =>
                           n9425, A => n28596, ZN => n28593);
   U21721 : OAI22_X1 port map( A1 => n9105, A2 => n30300, B1 => n9873, B2 => 
                           n30294, ZN => n28596);
   U21722 : AOI221_X1 port map( B1 => n30312, B2 => n22042, C1 => n30306, C2 =>
                           n9420, A => n28577, ZN => n28574);
   U21723 : OAI22_X1 port map( A1 => n9100, A2 => n30300, B1 => n9868, B2 => 
                           n30294, ZN => n28577);
   U21724 : AOI221_X1 port map( B1 => n30312, B2 => n22043, C1 => n30306, C2 =>
                           n9415, A => n28558, ZN => n28555);
   U21725 : OAI22_X1 port map( A1 => n9095, A2 => n30300, B1 => n9863, B2 => 
                           n30294, ZN => n28558);
   U21726 : AOI221_X1 port map( B1 => n30312, B2 => n22044, C1 => n30306, C2 =>
                           n9410, A => n28539, ZN => n28536);
   U21727 : OAI22_X1 port map( A1 => n9090, A2 => n30300, B1 => n9858, B2 => 
                           n30294, ZN => n28539);
   U21728 : AOI221_X1 port map( B1 => n30312, B2 => n22045, C1 => n30306, C2 =>
                           n9405, A => n28520, ZN => n28517);
   U21729 : OAI22_X1 port map( A1 => n9085, A2 => n30300, B1 => n9853, B2 => 
                           n30294, ZN => n28520);
   U21730 : AOI221_X1 port map( B1 => n30312, B2 => n22046, C1 => n30306, C2 =>
                           n9400, A => n28501, ZN => n28498);
   U21731 : OAI22_X1 port map( A1 => n9080, A2 => n30300, B1 => n9848, B2 => 
                           n30294, ZN => n28501);
   U21732 : AOI221_X1 port map( B1 => n30312, B2 => n22047, C1 => n30306, C2 =>
                           n9395, A => n28482, ZN => n28479);
   U21733 : OAI22_X1 port map( A1 => n9075, A2 => n30300, B1 => n9843, B2 => 
                           n30294, ZN => n28482);
   U21734 : AOI221_X1 port map( B1 => n30312, B2 => n22048, C1 => n30306, C2 =>
                           n9390, A => n28463, ZN => n28460);
   U21735 : OAI22_X1 port map( A1 => n9070, A2 => n30300, B1 => n9838, B2 => 
                           n30294, ZN => n28463);
   U21736 : AOI221_X1 port map( B1 => n30312, B2 => n22049, C1 => n30306, C2 =>
                           n9385, A => n28444, ZN => n28441);
   U21737 : OAI22_X1 port map( A1 => n9065, A2 => n30300, B1 => n9833, B2 => 
                           n30294, ZN => n28444);
   U21738 : AOI221_X1 port map( B1 => n30312, B2 => n22050, C1 => n30306, C2 =>
                           n9380, A => n28425, ZN => n28422);
   U21739 : OAI22_X1 port map( A1 => n9060, A2 => n30300, B1 => n9828, B2 => 
                           n30294, ZN => n28425);
   U21740 : AOI221_X1 port map( B1 => n30312, B2 => n22051, C1 => n30306, C2 =>
                           n9375, A => n28406, ZN => n28403);
   U21741 : OAI22_X1 port map( A1 => n9055, A2 => n30300, B1 => n9823, B2 => 
                           n30294, ZN => n28406);
   U21742 : AOI221_X1 port map( B1 => n30312, B2 => n22052, C1 => n30306, C2 =>
                           n9370, A => n28387, ZN => n28384);
   U21743 : OAI22_X1 port map( A1 => n9050, A2 => n30300, B1 => n9818, B2 => 
                           n30294, ZN => n28387);
   U21744 : AOI221_X1 port map( B1 => n30313, B2 => n22053, C1 => n30307, C2 =>
                           n9365, A => n28368, ZN => n28365);
   U21745 : OAI22_X1 port map( A1 => n9045, A2 => n30301, B1 => n9813, B2 => 
                           n30295, ZN => n28368);
   U21746 : AOI221_X1 port map( B1 => n30313, B2 => n22054, C1 => n30307, C2 =>
                           n9360, A => n28349, ZN => n28346);
   U21747 : OAI22_X1 port map( A1 => n9040, A2 => n30301, B1 => n9808, B2 => 
                           n30295, ZN => n28349);
   U21748 : AOI221_X1 port map( B1 => n30313, B2 => n22055, C1 => n30307, C2 =>
                           n9355, A => n28330, ZN => n28327);
   U21749 : OAI22_X1 port map( A1 => n9035, A2 => n30301, B1 => n9803, B2 => 
                           n30295, ZN => n28330);
   U21750 : AOI221_X1 port map( B1 => n30313, B2 => n22056, C1 => n30307, C2 =>
                           n9350, A => n28311, ZN => n28308);
   U21751 : OAI22_X1 port map( A1 => n9030, A2 => n30301, B1 => n9798, B2 => 
                           n30295, ZN => n28311);
   U21752 : AOI221_X1 port map( B1 => n30313, B2 => n22057, C1 => n30307, C2 =>
                           n9345, A => n28292, ZN => n28289);
   U21753 : OAI22_X1 port map( A1 => n9025, A2 => n30301, B1 => n9793, B2 => 
                           n30295, ZN => n28292);
   U21754 : AOI221_X1 port map( B1 => n30313, B2 => n22058, C1 => n30307, C2 =>
                           n9340, A => n28273, ZN => n28270);
   U21755 : OAI22_X1 port map( A1 => n9020, A2 => n30301, B1 => n9788, B2 => 
                           n30295, ZN => n28273);
   U21756 : AOI221_X1 port map( B1 => n30313, B2 => n22059, C1 => n30307, C2 =>
                           n9335, A => n28254, ZN => n28251);
   U21757 : OAI22_X1 port map( A1 => n9015, A2 => n30301, B1 => n9783, B2 => 
                           n30295, ZN => n28254);
   U21758 : AOI221_X1 port map( B1 => n30313, B2 => n22060, C1 => n30307, C2 =>
                           n9330, A => n28235, ZN => n28232);
   U21759 : OAI22_X1 port map( A1 => n9010, A2 => n30301, B1 => n9778, B2 => 
                           n30295, ZN => n28235);
   U21760 : AOI221_X1 port map( B1 => n30313, B2 => n22061, C1 => n30307, C2 =>
                           n9325, A => n28216, ZN => n28213);
   U21761 : OAI22_X1 port map( A1 => n9005, A2 => n30301, B1 => n9773, B2 => 
                           n30295, ZN => n28216);
   U21762 : AOI221_X1 port map( B1 => n30313, B2 => n22062, C1 => n30307, C2 =>
                           n9320, A => n28197, ZN => n28194);
   U21763 : OAI22_X1 port map( A1 => n9000, A2 => n30301, B1 => n9768, B2 => 
                           n30295, ZN => n28197);
   U21764 : AOI221_X1 port map( B1 => n30313, B2 => n22063, C1 => n30307, C2 =>
                           n9315, A => n28178, ZN => n28175);
   U21765 : OAI22_X1 port map( A1 => n8995, A2 => n30301, B1 => n9763, B2 => 
                           n30295, ZN => n28178);
   U21766 : AOI221_X1 port map( B1 => n30313, B2 => n22064, C1 => n30307, C2 =>
                           n9310, A => n28159, ZN => n28156);
   U21767 : OAI22_X1 port map( A1 => n8990, A2 => n30301, B1 => n9758, B2 => 
                           n30295, ZN => n28159);
   U21768 : AOI221_X1 port map( B1 => n30218, B2 => n21919, C1 => n30212, C2 =>
                           n9308, A => n28148, ZN => n28145);
   U21769 : OAI22_X1 port map( A1 => n26028, A2 => n30206, B1 => n25962, B2 => 
                           n30200, ZN => n28148);
   U21770 : AOI221_X1 port map( B1 => n30314, B2 => n21923, C1 => n30308, C2 =>
                           n9305, A => n28140, ZN => n28137);
   U21771 : OAI22_X1 port map( A1 => n8985, A2 => n30302, B1 => n9753, B2 => 
                           n30296, ZN => n28140);
   U21772 : AOI221_X1 port map( B1 => n30218, B2 => n21920, C1 => n30212, C2 =>
                           n9303, A => n28129, ZN => n28126);
   U21773 : OAI22_X1 port map( A1 => n26027, A2 => n30206, B1 => n25961, B2 => 
                           n30200, ZN => n28129);
   U21774 : AOI221_X1 port map( B1 => n30314, B2 => n21924, C1 => n30308, C2 =>
                           n9300, A => n28121, ZN => n28118);
   U21775 : OAI22_X1 port map( A1 => n8980, A2 => n30302, B1 => n9748, B2 => 
                           n30296, ZN => n28121);
   U21776 : AOI221_X1 port map( B1 => n30218, B2 => n21921, C1 => n30212, C2 =>
                           n9298, A => n28110, ZN => n28107);
   U21777 : OAI22_X1 port map( A1 => n26026, A2 => n30206, B1 => n25960, B2 => 
                           n30200, ZN => n28110);
   U21778 : AOI221_X1 port map( B1 => n30314, B2 => n21925, C1 => n30308, C2 =>
                           n9295, A => n28102, ZN => n28099);
   U21779 : OAI22_X1 port map( A1 => n8975, A2 => n30302, B1 => n9743, B2 => 
                           n30296, ZN => n28102);
   U21780 : AOI221_X1 port map( B1 => n30218, B2 => n21922, C1 => n30212, C2 =>
                           n9293, A => n28080, ZN => n28071);
   U21781 : OAI22_X1 port map( A1 => n26024, A2 => n30206, B1 => n25958, B2 => 
                           n30200, ZN => n28080);
   U21782 : AOI221_X1 port map( B1 => n30314, B2 => n21926, C1 => n30308, C2 =>
                           n9290, A => n28056, ZN => n28047);
   U21783 : OAI22_X1 port map( A1 => n8970, A2 => n30302, B1 => n9738, B2 => 
                           n30296, ZN => n28056);
   U21784 : AOI221_X1 port map( B1 => n30514, B2 => n22065, C1 => n30508, C2 =>
                           n9605, A => n28004, ZN => n27997);
   U21785 : OAI22_X1 port map( A1 => n9285, A2 => n30502, B1 => n25381, B2 => 
                           n30496, ZN => n28004);
   U21786 : AOI221_X1 port map( B1 => n30514, B2 => n22066, C1 => n30508, C2 =>
                           n9600, A => n27973, ZN => n27970);
   U21787 : OAI22_X1 port map( A1 => n9280, A2 => n30502, B1 => n25380, B2 => 
                           n30496, ZN => n27973);
   U21788 : AOI221_X1 port map( B1 => n30514, B2 => n22067, C1 => n30508, C2 =>
                           n9595, A => n27947, ZN => n27944);
   U21789 : OAI22_X1 port map( A1 => n9275, A2 => n30502, B1 => n25379, B2 => 
                           n30496, ZN => n27947);
   U21790 : AOI221_X1 port map( B1 => n30514, B2 => n22068, C1 => n30508, C2 =>
                           n9590, A => n27921, ZN => n27918);
   U21791 : OAI22_X1 port map( A1 => n9270, A2 => n30502, B1 => n25378, B2 => 
                           n30496, ZN => n27921);
   U21792 : AOI221_X1 port map( B1 => n30514, B2 => n22069, C1 => n30508, C2 =>
                           n9585, A => n27895, ZN => n27892);
   U21793 : OAI22_X1 port map( A1 => n9265, A2 => n30502, B1 => n25377, B2 => 
                           n30496, ZN => n27895);
   U21794 : AOI221_X1 port map( B1 => n30514, B2 => n22070, C1 => n30508, C2 =>
                           n9580, A => n27869, ZN => n27866);
   U21795 : OAI22_X1 port map( A1 => n9260, A2 => n30502, B1 => n25376, B2 => 
                           n30496, ZN => n27869);
   U21796 : AOI221_X1 port map( B1 => n30514, B2 => n22071, C1 => n30508, C2 =>
                           n9575, A => n27843, ZN => n27840);
   U21797 : OAI22_X1 port map( A1 => n9255, A2 => n30502, B1 => n25375, B2 => 
                           n30496, ZN => n27843);
   U21798 : AOI221_X1 port map( B1 => n30514, B2 => n22072, C1 => n30508, C2 =>
                           n9570, A => n27817, ZN => n27814);
   U21799 : OAI22_X1 port map( A1 => n9250, A2 => n30502, B1 => n25374, B2 => 
                           n30496, ZN => n27817);
   U21800 : AOI221_X1 port map( B1 => n30514, B2 => n22073, C1 => n30508, C2 =>
                           n9565, A => n27791, ZN => n27788);
   U21801 : OAI22_X1 port map( A1 => n9245, A2 => n30502, B1 => n25373, B2 => 
                           n30496, ZN => n27791);
   U21802 : AOI221_X1 port map( B1 => n30514, B2 => n22074, C1 => n30508, C2 =>
                           n9560, A => n27765, ZN => n27762);
   U21803 : OAI22_X1 port map( A1 => n9240, A2 => n30502, B1 => n25372, B2 => 
                           n30496, ZN => n27765);
   U21804 : AOI221_X1 port map( B1 => n30514, B2 => n22075, C1 => n30508, C2 =>
                           n9555, A => n27739, ZN => n27736);
   U21805 : OAI22_X1 port map( A1 => n9235, A2 => n30502, B1 => n25371, B2 => 
                           n30496, ZN => n27739);
   U21806 : AOI221_X1 port map( B1 => n30514, B2 => n22016, C1 => n30508, C2 =>
                           n9550, A => n27713, ZN => n27710);
   U21807 : OAI22_X1 port map( A1 => n9230, A2 => n30502, B1 => n9998, B2 => 
                           n30496, ZN => n27713);
   U21808 : AOI221_X1 port map( B1 => n30515, B2 => n22017, C1 => n30509, C2 =>
                           n9545, A => n27687, ZN => n27684);
   U21809 : OAI22_X1 port map( A1 => n9225, A2 => n30503, B1 => n9993, B2 => 
                           n30497, ZN => n27687);
   U21810 : AOI221_X1 port map( B1 => n30515, B2 => n22018, C1 => n30509, C2 =>
                           n9540, A => n27661, ZN => n27658);
   U21811 : OAI22_X1 port map( A1 => n9220, A2 => n30503, B1 => n9988, B2 => 
                           n30497, ZN => n27661);
   U21812 : AOI221_X1 port map( B1 => n30515, B2 => n22019, C1 => n30509, C2 =>
                           n9535, A => n27635, ZN => n27632);
   U21813 : OAI22_X1 port map( A1 => n9215, A2 => n30503, B1 => n9983, B2 => 
                           n30497, ZN => n27635);
   U21814 : AOI221_X1 port map( B1 => n30515, B2 => n22020, C1 => n30509, C2 =>
                           n9530, A => n27609, ZN => n27606);
   U21815 : OAI22_X1 port map( A1 => n9210, A2 => n30503, B1 => n9978, B2 => 
                           n30497, ZN => n27609);
   U21816 : AOI221_X1 port map( B1 => n30515, B2 => n22021, C1 => n30509, C2 =>
                           n9525, A => n27583, ZN => n27580);
   U21817 : OAI22_X1 port map( A1 => n9205, A2 => n30503, B1 => n9973, B2 => 
                           n30497, ZN => n27583);
   U21818 : AOI221_X1 port map( B1 => n30515, B2 => n22022, C1 => n30509, C2 =>
                           n9520, A => n27557, ZN => n27554);
   U21819 : OAI22_X1 port map( A1 => n9200, A2 => n30503, B1 => n9968, B2 => 
                           n30497, ZN => n27557);
   U21820 : AOI221_X1 port map( B1 => n30515, B2 => n22023, C1 => n30509, C2 =>
                           n9515, A => n27531, ZN => n27528);
   U21821 : OAI22_X1 port map( A1 => n9195, A2 => n30503, B1 => n9963, B2 => 
                           n30497, ZN => n27531);
   U21822 : AOI221_X1 port map( B1 => n30515, B2 => n22024, C1 => n30509, C2 =>
                           n9510, A => n27505, ZN => n27502);
   U21823 : OAI22_X1 port map( A1 => n9190, A2 => n30503, B1 => n9958, B2 => 
                           n30497, ZN => n27505);
   U21824 : AOI221_X1 port map( B1 => n30515, B2 => n22025, C1 => n30509, C2 =>
                           n9505, A => n27479, ZN => n27476);
   U21825 : OAI22_X1 port map( A1 => n9185, A2 => n30503, B1 => n9953, B2 => 
                           n30497, ZN => n27479);
   U21826 : AOI221_X1 port map( B1 => n30515, B2 => n22026, C1 => n30509, C2 =>
                           n9500, A => n27453, ZN => n27450);
   U21827 : OAI22_X1 port map( A1 => n9180, A2 => n30503, B1 => n9948, B2 => 
                           n30497, ZN => n27453);
   U21828 : AOI221_X1 port map( B1 => n30515, B2 => n22027, C1 => n30509, C2 =>
                           n9495, A => n27427, ZN => n27424);
   U21829 : OAI22_X1 port map( A1 => n9175, A2 => n30503, B1 => n9943, B2 => 
                           n30497, ZN => n27427);
   U21830 : AOI221_X1 port map( B1 => n30515, B2 => n22028, C1 => n30509, C2 =>
                           n9490, A => n27401, ZN => n27398);
   U21831 : OAI22_X1 port map( A1 => n9170, A2 => n30503, B1 => n9938, B2 => 
                           n30497, ZN => n27401);
   U21832 : AOI221_X1 port map( B1 => n30516, B2 => n22029, C1 => n30510, C2 =>
                           n9485, A => n27375, ZN => n27372);
   U21833 : OAI22_X1 port map( A1 => n9165, A2 => n30504, B1 => n9933, B2 => 
                           n30498, ZN => n27375);
   U21834 : AOI221_X1 port map( B1 => n30516, B2 => n22030, C1 => n30510, C2 =>
                           n9480, A => n27349, ZN => n27346);
   U21835 : OAI22_X1 port map( A1 => n9160, A2 => n30504, B1 => n9928, B2 => 
                           n30498, ZN => n27349);
   U21836 : AOI221_X1 port map( B1 => n30516, B2 => n22031, C1 => n30510, C2 =>
                           n9475, A => n27323, ZN => n27320);
   U21837 : OAI22_X1 port map( A1 => n9155, A2 => n30504, B1 => n9923, B2 => 
                           n30498, ZN => n27323);
   U21838 : AOI221_X1 port map( B1 => n30516, B2 => n22032, C1 => n30510, C2 =>
                           n9470, A => n27297, ZN => n27294);
   U21839 : OAI22_X1 port map( A1 => n9150, A2 => n30504, B1 => n9918, B2 => 
                           n30498, ZN => n27297);
   U21840 : AOI221_X1 port map( B1 => n30516, B2 => n22033, C1 => n30510, C2 =>
                           n9465, A => n27271, ZN => n27268);
   U21841 : OAI22_X1 port map( A1 => n9145, A2 => n30504, B1 => n9913, B2 => 
                           n30498, ZN => n27271);
   U21842 : AOI221_X1 port map( B1 => n30516, B2 => n22034, C1 => n30510, C2 =>
                           n9460, A => n27245, ZN => n27242);
   U21843 : OAI22_X1 port map( A1 => n9140, A2 => n30504, B1 => n9908, B2 => 
                           n30498, ZN => n27245);
   U21844 : AOI221_X1 port map( B1 => n30516, B2 => n22035, C1 => n30510, C2 =>
                           n9455, A => n27219, ZN => n27216);
   U21845 : OAI22_X1 port map( A1 => n9135, A2 => n30504, B1 => n9903, B2 => 
                           n30498, ZN => n27219);
   U21846 : AOI221_X1 port map( B1 => n30516, B2 => n22036, C1 => n30510, C2 =>
                           n9450, A => n27193, ZN => n27190);
   U21847 : OAI22_X1 port map( A1 => n9130, A2 => n30504, B1 => n9898, B2 => 
                           n30498, ZN => n27193);
   U21848 : AOI221_X1 port map( B1 => n30516, B2 => n22037, C1 => n30510, C2 =>
                           n9445, A => n27167, ZN => n27164);
   U21849 : OAI22_X1 port map( A1 => n9125, A2 => n30504, B1 => n9893, B2 => 
                           n30498, ZN => n27167);
   U21850 : AOI221_X1 port map( B1 => n30516, B2 => n22038, C1 => n30510, C2 =>
                           n9440, A => n27141, ZN => n27138);
   U21851 : OAI22_X1 port map( A1 => n9120, A2 => n30504, B1 => n9888, B2 => 
                           n30498, ZN => n27141);
   U21852 : AOI221_X1 port map( B1 => n30516, B2 => n22039, C1 => n30510, C2 =>
                           n9435, A => n27115, ZN => n27112);
   U21853 : OAI22_X1 port map( A1 => n9115, A2 => n30504, B1 => n9883, B2 => 
                           n30498, ZN => n27115);
   U21854 : AOI221_X1 port map( B1 => n30516, B2 => n22040, C1 => n30510, C2 =>
                           n9430, A => n27089, ZN => n27086);
   U21855 : OAI22_X1 port map( A1 => n9110, A2 => n30504, B1 => n9878, B2 => 
                           n30498, ZN => n27089);
   U21856 : AOI221_X1 port map( B1 => n30517, B2 => n22041, C1 => n30511, C2 =>
                           n9425, A => n27063, ZN => n27060);
   U21857 : OAI22_X1 port map( A1 => n9105, A2 => n30505, B1 => n9873, B2 => 
                           n30499, ZN => n27063);
   U21858 : AOI221_X1 port map( B1 => n30517, B2 => n22042, C1 => n30511, C2 =>
                           n9420, A => n27037, ZN => n27034);
   U21859 : OAI22_X1 port map( A1 => n9100, A2 => n30505, B1 => n9868, B2 => 
                           n30499, ZN => n27037);
   U21860 : AOI221_X1 port map( B1 => n30517, B2 => n22043, C1 => n30511, C2 =>
                           n9415, A => n27011, ZN => n27008);
   U21861 : OAI22_X1 port map( A1 => n9095, A2 => n30505, B1 => n9863, B2 => 
                           n30499, ZN => n27011);
   U21862 : AOI221_X1 port map( B1 => n30517, B2 => n22044, C1 => n30511, C2 =>
                           n9410, A => n26985, ZN => n26982);
   U21863 : OAI22_X1 port map( A1 => n9090, A2 => n30505, B1 => n9858, B2 => 
                           n30499, ZN => n26985);
   U21864 : AOI221_X1 port map( B1 => n30517, B2 => n22045, C1 => n30511, C2 =>
                           n9405, A => n26959, ZN => n26956);
   U21865 : OAI22_X1 port map( A1 => n9085, A2 => n30505, B1 => n9853, B2 => 
                           n30499, ZN => n26959);
   U21866 : AOI221_X1 port map( B1 => n30517, B2 => n22046, C1 => n30511, C2 =>
                           n9400, A => n26933, ZN => n26930);
   U21867 : OAI22_X1 port map( A1 => n9080, A2 => n30505, B1 => n9848, B2 => 
                           n30499, ZN => n26933);
   U21868 : AOI221_X1 port map( B1 => n30517, B2 => n22047, C1 => n30511, C2 =>
                           n9395, A => n26907, ZN => n26904);
   U21869 : OAI22_X1 port map( A1 => n9075, A2 => n30505, B1 => n9843, B2 => 
                           n30499, ZN => n26907);
   U21870 : AOI221_X1 port map( B1 => n30517, B2 => n22048, C1 => n30511, C2 =>
                           n9390, A => n26881, ZN => n26878);
   U21871 : OAI22_X1 port map( A1 => n9070, A2 => n30505, B1 => n9838, B2 => 
                           n30499, ZN => n26881);
   U21872 : AOI221_X1 port map( B1 => n30517, B2 => n22049, C1 => n30511, C2 =>
                           n9385, A => n26855, ZN => n26852);
   U21873 : OAI22_X1 port map( A1 => n9065, A2 => n30505, B1 => n9833, B2 => 
                           n30499, ZN => n26855);
   U21874 : AOI221_X1 port map( B1 => n30517, B2 => n22050, C1 => n30511, C2 =>
                           n9380, A => n26829, ZN => n26826);
   U21875 : OAI22_X1 port map( A1 => n9060, A2 => n30505, B1 => n9828, B2 => 
                           n30499, ZN => n26829);
   U21876 : AOI221_X1 port map( B1 => n30517, B2 => n22051, C1 => n30511, C2 =>
                           n9375, A => n26803, ZN => n26800);
   U21877 : OAI22_X1 port map( A1 => n9055, A2 => n30505, B1 => n9823, B2 => 
                           n30499, ZN => n26803);
   U21878 : AOI221_X1 port map( B1 => n30517, B2 => n22052, C1 => n30511, C2 =>
                           n9370, A => n26777, ZN => n26774);
   U21879 : OAI22_X1 port map( A1 => n9050, A2 => n30505, B1 => n9818, B2 => 
                           n30499, ZN => n26777);
   U21880 : AOI221_X1 port map( B1 => n30518, B2 => n22053, C1 => n30512, C2 =>
                           n9365, A => n26751, ZN => n26748);
   U21881 : OAI22_X1 port map( A1 => n9045, A2 => n30506, B1 => n9813, B2 => 
                           n30500, ZN => n26751);
   U21882 : AOI221_X1 port map( B1 => n30518, B2 => n22054, C1 => n30512, C2 =>
                           n9360, A => n26725, ZN => n26722);
   U21883 : OAI22_X1 port map( A1 => n9040, A2 => n30506, B1 => n9808, B2 => 
                           n30500, ZN => n26725);
   U21884 : AOI221_X1 port map( B1 => n30518, B2 => n22055, C1 => n30512, C2 =>
                           n9355, A => n26699, ZN => n26696);
   U21885 : OAI22_X1 port map( A1 => n9035, A2 => n30506, B1 => n9803, B2 => 
                           n30500, ZN => n26699);
   U21886 : AOI221_X1 port map( B1 => n30518, B2 => n22056, C1 => n30512, C2 =>
                           n9350, A => n26673, ZN => n26670);
   U21887 : OAI22_X1 port map( A1 => n9030, A2 => n30506, B1 => n9798, B2 => 
                           n30500, ZN => n26673);
   U21888 : AOI221_X1 port map( B1 => n30518, B2 => n22057, C1 => n30512, C2 =>
                           n9345, A => n26647, ZN => n26644);
   U21889 : OAI22_X1 port map( A1 => n9025, A2 => n30506, B1 => n9793, B2 => 
                           n30500, ZN => n26647);
   U21890 : AOI221_X1 port map( B1 => n30518, B2 => n22058, C1 => n30512, C2 =>
                           n9340, A => n26621, ZN => n26618);
   U21891 : OAI22_X1 port map( A1 => n9020, A2 => n30506, B1 => n9788, B2 => 
                           n30500, ZN => n26621);
   U21892 : AOI221_X1 port map( B1 => n30518, B2 => n22059, C1 => n30512, C2 =>
                           n9335, A => n26595, ZN => n26592);
   U21893 : OAI22_X1 port map( A1 => n9015, A2 => n30506, B1 => n9783, B2 => 
                           n30500, ZN => n26595);
   U21894 : AOI221_X1 port map( B1 => n30518, B2 => n22060, C1 => n30512, C2 =>
                           n9330, A => n26569, ZN => n26566);
   U21895 : OAI22_X1 port map( A1 => n9010, A2 => n30506, B1 => n9778, B2 => 
                           n30500, ZN => n26569);
   U21896 : AOI221_X1 port map( B1 => n30518, B2 => n22061, C1 => n30512, C2 =>
                           n9325, A => n26543, ZN => n26540);
   U21897 : OAI22_X1 port map( A1 => n9005, A2 => n30506, B1 => n9773, B2 => 
                           n30500, ZN => n26543);
   U21898 : AOI221_X1 port map( B1 => n30518, B2 => n22062, C1 => n30512, C2 =>
                           n9320, A => n26517, ZN => n26514);
   U21899 : OAI22_X1 port map( A1 => n9000, A2 => n30506, B1 => n9768, B2 => 
                           n30500, ZN => n26517);
   U21900 : AOI221_X1 port map( B1 => n30518, B2 => n22063, C1 => n30512, C2 =>
                           n9315, A => n26491, ZN => n26488);
   U21901 : OAI22_X1 port map( A1 => n8995, A2 => n30506, B1 => n9763, B2 => 
                           n30500, ZN => n26491);
   U21902 : AOI221_X1 port map( B1 => n30518, B2 => n22064, C1 => n30512, C2 =>
                           n9310, A => n26465, ZN => n26462);
   U21903 : OAI22_X1 port map( A1 => n8990, A2 => n30506, B1 => n9758, B2 => 
                           n30500, ZN => n26465);
   U21904 : AOI221_X1 port map( B1 => n30519, B2 => n21923, C1 => n30513, C2 =>
                           n9305, A => n26439, ZN => n26436);
   U21905 : OAI22_X1 port map( A1 => n8985, A2 => n30507, B1 => n9753, B2 => 
                           n30501, ZN => n26439);
   U21906 : AOI221_X1 port map( B1 => n30519, B2 => n21924, C1 => n30513, C2 =>
                           n9300, A => n26413, ZN => n26410);
   U21907 : OAI22_X1 port map( A1 => n8980, A2 => n30507, B1 => n9748, B2 => 
                           n30501, ZN => n26413);
   U21908 : AOI221_X1 port map( B1 => n30519, B2 => n21925, C1 => n30513, C2 =>
                           n9295, A => n26387, ZN => n26384);
   U21909 : OAI22_X1 port map( A1 => n8975, A2 => n30507, B1 => n9743, B2 => 
                           n30501, ZN => n26387);
   U21910 : AOI221_X1 port map( B1 => n30519, B2 => n21926, C1 => n30513, C2 =>
                           n9290, A => n26335, ZN => n26326);
   U21911 : OAI22_X1 port map( A1 => n8970, A2 => n30507, B1 => n9738, B2 => 
                           n30501, ZN => n26335);
   U21912 : AOI221_X1 port map( B1 => n30417, B2 => n29764, C1 => n30411, C2 =>
                           n29572, A => n28023, ZN => n28016);
   U21913 : OAI22_X1 port map( A1 => n9286, A2 => n30405, B1 => n25667, B2 => 
                           n30399, ZN => n28023);
   U21914 : AOI221_X1 port map( B1 => n30417, B2 => n29765, C1 => n30411, C2 =>
                           n29573, A => n27983, ZN => n27978);
   U21915 : OAI22_X1 port map( A1 => n9281, A2 => n30405, B1 => n25666, B2 => 
                           n30399, ZN => n27983);
   U21916 : AOI221_X1 port map( B1 => n30417, B2 => n29766, C1 => n30411, C2 =>
                           n29574, A => n27957, ZN => n27952);
   U21917 : OAI22_X1 port map( A1 => n9276, A2 => n30405, B1 => n25665, B2 => 
                           n30399, ZN => n27957);
   U21918 : AOI221_X1 port map( B1 => n30417, B2 => n29767, C1 => n30411, C2 =>
                           n29575, A => n27931, ZN => n27926);
   U21919 : OAI22_X1 port map( A1 => n9271, A2 => n30405, B1 => n25664, B2 => 
                           n30399, ZN => n27931);
   U21920 : AOI221_X1 port map( B1 => n30417, B2 => n29768, C1 => n30411, C2 =>
                           n29576, A => n27905, ZN => n27900);
   U21921 : OAI22_X1 port map( A1 => n9266, A2 => n30405, B1 => n25663, B2 => 
                           n30399, ZN => n27905);
   U21922 : AOI221_X1 port map( B1 => n30417, B2 => n29769, C1 => n30411, C2 =>
                           n29577, A => n27879, ZN => n27874);
   U21923 : OAI22_X1 port map( A1 => n9261, A2 => n30405, B1 => n25662, B2 => 
                           n30399, ZN => n27879);
   U21924 : AOI221_X1 port map( B1 => n30417, B2 => n29770, C1 => n30411, C2 =>
                           n29578, A => n27853, ZN => n27848);
   U21925 : OAI22_X1 port map( A1 => n9256, A2 => n30405, B1 => n25661, B2 => 
                           n30399, ZN => n27853);
   U21926 : AOI221_X1 port map( B1 => n30417, B2 => n29771, C1 => n30411, C2 =>
                           n29579, A => n27827, ZN => n27822);
   U21927 : OAI22_X1 port map( A1 => n9251, A2 => n30405, B1 => n25660, B2 => 
                           n30399, ZN => n27827);
   U21928 : AOI221_X1 port map( B1 => n30417, B2 => n29772, C1 => n30411, C2 =>
                           n29580, A => n27801, ZN => n27796);
   U21929 : OAI22_X1 port map( A1 => n9246, A2 => n30405, B1 => n25659, B2 => 
                           n30399, ZN => n27801);
   U21930 : AOI221_X1 port map( B1 => n30417, B2 => n29773, C1 => n30411, C2 =>
                           n29581, A => n27775, ZN => n27770);
   U21931 : OAI22_X1 port map( A1 => n9241, A2 => n30405, B1 => n25658, B2 => 
                           n30399, ZN => n27775);
   U21932 : AOI221_X1 port map( B1 => n30417, B2 => n29774, C1 => n30411, C2 =>
                           n29582, A => n27749, ZN => n27744);
   U21933 : OAI22_X1 port map( A1 => n9236, A2 => n30405, B1 => n25657, B2 => 
                           n30399, ZN => n27749);
   U21934 : AOI221_X1 port map( B1 => n30417, B2 => n29775, C1 => n30411, C2 =>
                           n29583, A => n27723, ZN => n27718);
   U21935 : OAI22_X1 port map( A1 => n9231, A2 => n30405, B1 => n9999, B2 => 
                           n30399, ZN => n27723);
   U21936 : AOI221_X1 port map( B1 => n30418, B2 => n29776, C1 => n30412, C2 =>
                           n29584, A => n27697, ZN => n27692);
   U21937 : OAI22_X1 port map( A1 => n9226, A2 => n30406, B1 => n9994, B2 => 
                           n30400, ZN => n27697);
   U21938 : AOI221_X1 port map( B1 => n30418, B2 => n29777, C1 => n30412, C2 =>
                           n29585, A => n27671, ZN => n27666);
   U21939 : OAI22_X1 port map( A1 => n9221, A2 => n30406, B1 => n9989, B2 => 
                           n30400, ZN => n27671);
   U21940 : AOI221_X1 port map( B1 => n30418, B2 => n29778, C1 => n30412, C2 =>
                           n29586, A => n27645, ZN => n27640);
   U21941 : OAI22_X1 port map( A1 => n9216, A2 => n30406, B1 => n9984, B2 => 
                           n30400, ZN => n27645);
   U21942 : AOI221_X1 port map( B1 => n30418, B2 => n29779, C1 => n30412, C2 =>
                           n29587, A => n27619, ZN => n27614);
   U21943 : OAI22_X1 port map( A1 => n9211, A2 => n30406, B1 => n9979, B2 => 
                           n30400, ZN => n27619);
   U21944 : AOI221_X1 port map( B1 => n30418, B2 => n29780, C1 => n30412, C2 =>
                           n29588, A => n27593, ZN => n27588);
   U21945 : OAI22_X1 port map( A1 => n9206, A2 => n30406, B1 => n9974, B2 => 
                           n30400, ZN => n27593);
   U21946 : AOI221_X1 port map( B1 => n30418, B2 => n29781, C1 => n30412, C2 =>
                           n29589, A => n27567, ZN => n27562);
   U21947 : OAI22_X1 port map( A1 => n9201, A2 => n30406, B1 => n9969, B2 => 
                           n30400, ZN => n27567);
   U21948 : AOI221_X1 port map( B1 => n30418, B2 => n29782, C1 => n30412, C2 =>
                           n29590, A => n27541, ZN => n27536);
   U21949 : OAI22_X1 port map( A1 => n9196, A2 => n30406, B1 => n9964, B2 => 
                           n30400, ZN => n27541);
   U21950 : AOI221_X1 port map( B1 => n30418, B2 => n29783, C1 => n30412, C2 =>
                           n29591, A => n27515, ZN => n27510);
   U21951 : OAI22_X1 port map( A1 => n9191, A2 => n30406, B1 => n9959, B2 => 
                           n30400, ZN => n27515);
   U21952 : AOI221_X1 port map( B1 => n30418, B2 => n29784, C1 => n30412, C2 =>
                           n29592, A => n27489, ZN => n27484);
   U21953 : OAI22_X1 port map( A1 => n9186, A2 => n30406, B1 => n9954, B2 => 
                           n30400, ZN => n27489);
   U21954 : AOI221_X1 port map( B1 => n30418, B2 => n29785, C1 => n30412, C2 =>
                           n29593, A => n27463, ZN => n27458);
   U21955 : OAI22_X1 port map( A1 => n9181, A2 => n30406, B1 => n9949, B2 => 
                           n30400, ZN => n27463);
   U21956 : AOI221_X1 port map( B1 => n30418, B2 => n29786, C1 => n30412, C2 =>
                           n29594, A => n27437, ZN => n27432);
   U21957 : OAI22_X1 port map( A1 => n9176, A2 => n30406, B1 => n9944, B2 => 
                           n30400, ZN => n27437);
   U21958 : AOI221_X1 port map( B1 => n30418, B2 => n29787, C1 => n30412, C2 =>
                           n29595, A => n27411, ZN => n27406);
   U21959 : OAI22_X1 port map( A1 => n9171, A2 => n30406, B1 => n9939, B2 => 
                           n30400, ZN => n27411);
   U21960 : AOI221_X1 port map( B1 => n30419, B2 => n29788, C1 => n30413, C2 =>
                           n29596, A => n27385, ZN => n27380);
   U21961 : OAI22_X1 port map( A1 => n9166, A2 => n30407, B1 => n9934, B2 => 
                           n30401, ZN => n27385);
   U21962 : AOI221_X1 port map( B1 => n30419, B2 => n29789, C1 => n30413, C2 =>
                           n29597, A => n27359, ZN => n27354);
   U21963 : OAI22_X1 port map( A1 => n9161, A2 => n30407, B1 => n9929, B2 => 
                           n30401, ZN => n27359);
   U21964 : AOI221_X1 port map( B1 => n30419, B2 => n29790, C1 => n30413, C2 =>
                           n29598, A => n27333, ZN => n27328);
   U21965 : OAI22_X1 port map( A1 => n9156, A2 => n30407, B1 => n9924, B2 => 
                           n30401, ZN => n27333);
   U21966 : AOI221_X1 port map( B1 => n30419, B2 => n29791, C1 => n30413, C2 =>
                           n29599, A => n27307, ZN => n27302);
   U21967 : OAI22_X1 port map( A1 => n9151, A2 => n30407, B1 => n9919, B2 => 
                           n30401, ZN => n27307);
   U21968 : AOI221_X1 port map( B1 => n30419, B2 => n29792, C1 => n30413, C2 =>
                           n29600, A => n27281, ZN => n27276);
   U21969 : OAI22_X1 port map( A1 => n9146, A2 => n30407, B1 => n9914, B2 => 
                           n30401, ZN => n27281);
   U21970 : AOI221_X1 port map( B1 => n30419, B2 => n29793, C1 => n30413, C2 =>
                           n29601, A => n27255, ZN => n27250);
   U21971 : OAI22_X1 port map( A1 => n9141, A2 => n30407, B1 => n9909, B2 => 
                           n30401, ZN => n27255);
   U21972 : AOI221_X1 port map( B1 => n30419, B2 => n29794, C1 => n30413, C2 =>
                           n29602, A => n27229, ZN => n27224);
   U21973 : OAI22_X1 port map( A1 => n9136, A2 => n30407, B1 => n9904, B2 => 
                           n30401, ZN => n27229);
   U21974 : AOI221_X1 port map( B1 => n30419, B2 => n29795, C1 => n30413, C2 =>
                           n29603, A => n27203, ZN => n27198);
   U21975 : OAI22_X1 port map( A1 => n9131, A2 => n30407, B1 => n9899, B2 => 
                           n30401, ZN => n27203);
   U21976 : AOI221_X1 port map( B1 => n30419, B2 => n29796, C1 => n30413, C2 =>
                           n29604, A => n27177, ZN => n27172);
   U21977 : OAI22_X1 port map( A1 => n9126, A2 => n30407, B1 => n9894, B2 => 
                           n30401, ZN => n27177);
   U21978 : AOI221_X1 port map( B1 => n30419, B2 => n29797, C1 => n30413, C2 =>
                           n29605, A => n27151, ZN => n27146);
   U21979 : OAI22_X1 port map( A1 => n9121, A2 => n30407, B1 => n9889, B2 => 
                           n30401, ZN => n27151);
   U21980 : AOI221_X1 port map( B1 => n30419, B2 => n29798, C1 => n30413, C2 =>
                           n29606, A => n27125, ZN => n27120);
   U21981 : OAI22_X1 port map( A1 => n9116, A2 => n30407, B1 => n9884, B2 => 
                           n30401, ZN => n27125);
   U21982 : AOI221_X1 port map( B1 => n30419, B2 => n29799, C1 => n30413, C2 =>
                           n29607, A => n27099, ZN => n27094);
   U21983 : OAI22_X1 port map( A1 => n9111, A2 => n30407, B1 => n9879, B2 => 
                           n30401, ZN => n27099);
   U21984 : AOI221_X1 port map( B1 => n30420, B2 => n29800, C1 => n30414, C2 =>
                           n29608, A => n27073, ZN => n27068);
   U21985 : OAI22_X1 port map( A1 => n9106, A2 => n30408, B1 => n9874, B2 => 
                           n30402, ZN => n27073);
   U21986 : AOI221_X1 port map( B1 => n30420, B2 => n29801, C1 => n30414, C2 =>
                           n29609, A => n27047, ZN => n27042);
   U21987 : OAI22_X1 port map( A1 => n9101, A2 => n30408, B1 => n9869, B2 => 
                           n30402, ZN => n27047);
   U21988 : AOI221_X1 port map( B1 => n30420, B2 => n29802, C1 => n30414, C2 =>
                           n29610, A => n27021, ZN => n27016);
   U21989 : OAI22_X1 port map( A1 => n9096, A2 => n30408, B1 => n9864, B2 => 
                           n30402, ZN => n27021);
   U21990 : AOI221_X1 port map( B1 => n30420, B2 => n29803, C1 => n30414, C2 =>
                           n29611, A => n26995, ZN => n26990);
   U21991 : OAI22_X1 port map( A1 => n9091, A2 => n30408, B1 => n9859, B2 => 
                           n30402, ZN => n26995);
   U21992 : AOI221_X1 port map( B1 => n30420, B2 => n29804, C1 => n30414, C2 =>
                           n29612, A => n26969, ZN => n26964);
   U21993 : OAI22_X1 port map( A1 => n9086, A2 => n30408, B1 => n9854, B2 => 
                           n30402, ZN => n26969);
   U21994 : AOI221_X1 port map( B1 => n30420, B2 => n29805, C1 => n30414, C2 =>
                           n29613, A => n26943, ZN => n26938);
   U21995 : OAI22_X1 port map( A1 => n9081, A2 => n30408, B1 => n9849, B2 => 
                           n30402, ZN => n26943);
   U21996 : AOI221_X1 port map( B1 => n30420, B2 => n29806, C1 => n30414, C2 =>
                           n29614, A => n26917, ZN => n26912);
   U21997 : OAI22_X1 port map( A1 => n9076, A2 => n30408, B1 => n9844, B2 => 
                           n30402, ZN => n26917);
   U21998 : AOI221_X1 port map( B1 => n30420, B2 => n29807, C1 => n30414, C2 =>
                           n29615, A => n26891, ZN => n26886);
   U21999 : OAI22_X1 port map( A1 => n9071, A2 => n30408, B1 => n9839, B2 => 
                           n30402, ZN => n26891);
   U22000 : AOI221_X1 port map( B1 => n30420, B2 => n29808, C1 => n30414, C2 =>
                           n29616, A => n26865, ZN => n26860);
   U22001 : OAI22_X1 port map( A1 => n9066, A2 => n30408, B1 => n9834, B2 => 
                           n30402, ZN => n26865);
   U22002 : AOI221_X1 port map( B1 => n30420, B2 => n29809, C1 => n30414, C2 =>
                           n29617, A => n26839, ZN => n26834);
   U22003 : OAI22_X1 port map( A1 => n9061, A2 => n30408, B1 => n9829, B2 => 
                           n30402, ZN => n26839);
   U22004 : AOI221_X1 port map( B1 => n30420, B2 => n29810, C1 => n30414, C2 =>
                           n29618, A => n26813, ZN => n26808);
   U22005 : OAI22_X1 port map( A1 => n9056, A2 => n30408, B1 => n9824, B2 => 
                           n30402, ZN => n26813);
   U22006 : AOI221_X1 port map( B1 => n30420, B2 => n29811, C1 => n30414, C2 =>
                           n29619, A => n26787, ZN => n26782);
   U22007 : OAI22_X1 port map( A1 => n9051, A2 => n30408, B1 => n9819, B2 => 
                           n30402, ZN => n26787);
   U22008 : AOI221_X1 port map( B1 => n30421, B2 => n29812, C1 => n30415, C2 =>
                           n29620, A => n26761, ZN => n26756);
   U22009 : OAI22_X1 port map( A1 => n9046, A2 => n30409, B1 => n9814, B2 => 
                           n30403, ZN => n26761);
   U22010 : AOI221_X1 port map( B1 => n30421, B2 => n29813, C1 => n30415, C2 =>
                           n29621, A => n26735, ZN => n26730);
   U22011 : OAI22_X1 port map( A1 => n9041, A2 => n30409, B1 => n9809, B2 => 
                           n30403, ZN => n26735);
   U22012 : AOI221_X1 port map( B1 => n30421, B2 => n29814, C1 => n30415, C2 =>
                           n29622, A => n26709, ZN => n26704);
   U22013 : OAI22_X1 port map( A1 => n9036, A2 => n30409, B1 => n9804, B2 => 
                           n30403, ZN => n26709);
   U22014 : AOI221_X1 port map( B1 => n30421, B2 => n29815, C1 => n30415, C2 =>
                           n29623, A => n26683, ZN => n26678);
   U22015 : OAI22_X1 port map( A1 => n9031, A2 => n30409, B1 => n9799, B2 => 
                           n30403, ZN => n26683);
   U22016 : AOI221_X1 port map( B1 => n30421, B2 => n29816, C1 => n30415, C2 =>
                           n29624, A => n26657, ZN => n26652);
   U22017 : OAI22_X1 port map( A1 => n9026, A2 => n30409, B1 => n9794, B2 => 
                           n30403, ZN => n26657);
   U22018 : AOI221_X1 port map( B1 => n30421, B2 => n29817, C1 => n30415, C2 =>
                           n29625, A => n26631, ZN => n26626);
   U22019 : OAI22_X1 port map( A1 => n9021, A2 => n30409, B1 => n9789, B2 => 
                           n30403, ZN => n26631);
   U22020 : AOI221_X1 port map( B1 => n30421, B2 => n29818, C1 => n30415, C2 =>
                           n29626, A => n26605, ZN => n26600);
   U22021 : OAI22_X1 port map( A1 => n9016, A2 => n30409, B1 => n9784, B2 => 
                           n30403, ZN => n26605);
   U22022 : AOI221_X1 port map( B1 => n30421, B2 => n29819, C1 => n30415, C2 =>
                           n29627, A => n26579, ZN => n26574);
   U22023 : OAI22_X1 port map( A1 => n9011, A2 => n30409, B1 => n9779, B2 => 
                           n30403, ZN => n26579);
   U22024 : AOI221_X1 port map( B1 => n30421, B2 => n29820, C1 => n30415, C2 =>
                           n29628, A => n26553, ZN => n26548);
   U22025 : OAI22_X1 port map( A1 => n9006, A2 => n30409, B1 => n9774, B2 => 
                           n30403, ZN => n26553);
   U22026 : AOI221_X1 port map( B1 => n30421, B2 => n29821, C1 => n30415, C2 =>
                           n29629, A => n26527, ZN => n26522);
   U22027 : OAI22_X1 port map( A1 => n9001, A2 => n30409, B1 => n9769, B2 => 
                           n30403, ZN => n26527);
   U22028 : AOI221_X1 port map( B1 => n30421, B2 => n29822, C1 => n30415, C2 =>
                           n29630, A => n26501, ZN => n26496);
   U22029 : OAI22_X1 port map( A1 => n8996, A2 => n30409, B1 => n9764, B2 => 
                           n30403, ZN => n26501);
   U22030 : AOI221_X1 port map( B1 => n30421, B2 => n29823, C1 => n30415, C2 =>
                           n29631, A => n26475, ZN => n26470);
   U22031 : OAI22_X1 port map( A1 => n8991, A2 => n30409, B1 => n9759, B2 => 
                           n30403, ZN => n26475);
   U22032 : AOI221_X1 port map( B1 => n30422, B2 => n29824, C1 => n30416, C2 =>
                           n29632, A => n26449, ZN => n26444);
   U22033 : OAI22_X1 port map( A1 => n8986, A2 => n30410, B1 => n9754, B2 => 
                           n30404, ZN => n26449);
   U22034 : AOI221_X1 port map( B1 => n30422, B2 => n29825, C1 => n30416, C2 =>
                           n29633, A => n26423, ZN => n26418);
   U22035 : OAI22_X1 port map( A1 => n8981, A2 => n30410, B1 => n9749, B2 => 
                           n30404, ZN => n26423);
   U22036 : AOI221_X1 port map( B1 => n30422, B2 => n29826, C1 => n30416, C2 =>
                           n29634, A => n26397, ZN => n26392);
   U22037 : OAI22_X1 port map( A1 => n8976, A2 => n30410, B1 => n9744, B2 => 
                           n30404, ZN => n26397);
   U22038 : AOI221_X1 port map( B1 => n30422, B2 => n29827, C1 => n30416, C2 =>
                           n29635, A => n26361, ZN => n26350);
   U22039 : OAI22_X1 port map( A1 => n8971, A2 => n30410, B1 => n9739, B2 => 
                           n30404, ZN => n26361);
   U22040 : AOI221_X1 port map( B1 => n30490, B2 => n21927, C1 => n30484, C2 =>
                           n9606, A => n28008, ZN => n27996);
   U22041 : OAI22_X1 port map( A1 => n25801, A2 => n30478, B1 => n25735, B2 => 
                           n30472, ZN => n28008);
   U22042 : AOI221_X1 port map( B1 => n30490, B2 => n21928, C1 => n30484, C2 =>
                           n9601, A => n27974, ZN => n27969);
   U22043 : OAI22_X1 port map( A1 => n25800, A2 => n30478, B1 => n25734, B2 => 
                           n30472, ZN => n27974);
   U22044 : AOI221_X1 port map( B1 => n30490, B2 => n21929, C1 => n30484, C2 =>
                           n9596, A => n27948, ZN => n27943);
   U22045 : OAI22_X1 port map( A1 => n25799, A2 => n30478, B1 => n25733, B2 => 
                           n30472, ZN => n27948);
   U22046 : AOI221_X1 port map( B1 => n30490, B2 => n21930, C1 => n30484, C2 =>
                           n9591, A => n27922, ZN => n27917);
   U22047 : OAI22_X1 port map( A1 => n25798, A2 => n30478, B1 => n25732, B2 => 
                           n30472, ZN => n27922);
   U22048 : AOI221_X1 port map( B1 => n30490, B2 => n21931, C1 => n30484, C2 =>
                           n9586, A => n27896, ZN => n27891);
   U22049 : OAI22_X1 port map( A1 => n25797, A2 => n30478, B1 => n25731, B2 => 
                           n30472, ZN => n27896);
   U22050 : AOI221_X1 port map( B1 => n30490, B2 => n21932, C1 => n30484, C2 =>
                           n9581, A => n27870, ZN => n27865);
   U22051 : OAI22_X1 port map( A1 => n25796, A2 => n30478, B1 => n25730, B2 => 
                           n30472, ZN => n27870);
   U22052 : AOI221_X1 port map( B1 => n30490, B2 => n21933, C1 => n30484, C2 =>
                           n9576, A => n27844, ZN => n27839);
   U22053 : OAI22_X1 port map( A1 => n25795, A2 => n30478, B1 => n25729, B2 => 
                           n30472, ZN => n27844);
   U22054 : AOI221_X1 port map( B1 => n30490, B2 => n21934, C1 => n30484, C2 =>
                           n9571, A => n27818, ZN => n27813);
   U22055 : OAI22_X1 port map( A1 => n25794, A2 => n30478, B1 => n25728, B2 => 
                           n30472, ZN => n27818);
   U22056 : AOI221_X1 port map( B1 => n30490, B2 => n21935, C1 => n30484, C2 =>
                           n9566, A => n27792, ZN => n27787);
   U22057 : OAI22_X1 port map( A1 => n25793, A2 => n30478, B1 => n25727, B2 => 
                           n30472, ZN => n27792);
   U22058 : AOI221_X1 port map( B1 => n30490, B2 => n21936, C1 => n30484, C2 =>
                           n9561, A => n27766, ZN => n27761);
   U22059 : OAI22_X1 port map( A1 => n25792, A2 => n30478, B1 => n25726, B2 => 
                           n30472, ZN => n27766);
   U22060 : AOI221_X1 port map( B1 => n30490, B2 => n21937, C1 => n30484, C2 =>
                           n9556, A => n27740, ZN => n27735);
   U22061 : OAI22_X1 port map( A1 => n25791, A2 => n30478, B1 => n25725, B2 => 
                           n30472, ZN => n27740);
   U22062 : AOI221_X1 port map( B1 => n30490, B2 => n21938, C1 => n30484, C2 =>
                           n9551, A => n27714, ZN => n27709);
   U22063 : OAI22_X1 port map( A1 => n25790, A2 => n30478, B1 => n25724, B2 => 
                           n30472, ZN => n27714);
   U22064 : AOI221_X1 port map( B1 => n30491, B2 => n21939, C1 => n30485, C2 =>
                           n9546, A => n27688, ZN => n27683);
   U22065 : OAI22_X1 port map( A1 => n25789, A2 => n30479, B1 => n25723, B2 => 
                           n30473, ZN => n27688);
   U22066 : AOI221_X1 port map( B1 => n30491, B2 => n21940, C1 => n30485, C2 =>
                           n9541, A => n27662, ZN => n27657);
   U22067 : OAI22_X1 port map( A1 => n25788, A2 => n30479, B1 => n25722, B2 => 
                           n30473, ZN => n27662);
   U22068 : AOI221_X1 port map( B1 => n30491, B2 => n21941, C1 => n30485, C2 =>
                           n9536, A => n27636, ZN => n27631);
   U22069 : OAI22_X1 port map( A1 => n25787, A2 => n30479, B1 => n25721, B2 => 
                           n30473, ZN => n27636);
   U22070 : AOI221_X1 port map( B1 => n30491, B2 => n21942, C1 => n30485, C2 =>
                           n9531, A => n27610, ZN => n27605);
   U22071 : OAI22_X1 port map( A1 => n25786, A2 => n30479, B1 => n25720, B2 => 
                           n30473, ZN => n27610);
   U22072 : AOI221_X1 port map( B1 => n30491, B2 => n21943, C1 => n30485, C2 =>
                           n9526, A => n27584, ZN => n27579);
   U22073 : OAI22_X1 port map( A1 => n25785, A2 => n30479, B1 => n25719, B2 => 
                           n30473, ZN => n27584);
   U22074 : AOI221_X1 port map( B1 => n30491, B2 => n21944, C1 => n30485, C2 =>
                           n9521, A => n27558, ZN => n27553);
   U22075 : OAI22_X1 port map( A1 => n25784, A2 => n30479, B1 => n25718, B2 => 
                           n30473, ZN => n27558);
   U22076 : AOI221_X1 port map( B1 => n30491, B2 => n21945, C1 => n30485, C2 =>
                           n9516, A => n27532, ZN => n27527);
   U22077 : OAI22_X1 port map( A1 => n25783, A2 => n30479, B1 => n25717, B2 => 
                           n30473, ZN => n27532);
   U22078 : AOI221_X1 port map( B1 => n30491, B2 => n21946, C1 => n30485, C2 =>
                           n9511, A => n27506, ZN => n27501);
   U22079 : OAI22_X1 port map( A1 => n25782, A2 => n30479, B1 => n25716, B2 => 
                           n30473, ZN => n27506);
   U22080 : AOI221_X1 port map( B1 => n30491, B2 => n21947, C1 => n30485, C2 =>
                           n9506, A => n27480, ZN => n27475);
   U22081 : OAI22_X1 port map( A1 => n25781, A2 => n30479, B1 => n25715, B2 => 
                           n30473, ZN => n27480);
   U22082 : AOI221_X1 port map( B1 => n30491, B2 => n21948, C1 => n30485, C2 =>
                           n9501, A => n27454, ZN => n27449);
   U22083 : OAI22_X1 port map( A1 => n25780, A2 => n30479, B1 => n25714, B2 => 
                           n30473, ZN => n27454);
   U22084 : AOI221_X1 port map( B1 => n30491, B2 => n21949, C1 => n30485, C2 =>
                           n9496, A => n27428, ZN => n27423);
   U22085 : OAI22_X1 port map( A1 => n25779, A2 => n30479, B1 => n25713, B2 => 
                           n30473, ZN => n27428);
   U22086 : AOI221_X1 port map( B1 => n30491, B2 => n21950, C1 => n30485, C2 =>
                           n9491, A => n27402, ZN => n27397);
   U22087 : OAI22_X1 port map( A1 => n25778, A2 => n30479, B1 => n25712, B2 => 
                           n30473, ZN => n27402);
   U22088 : AOI221_X1 port map( B1 => n30492, B2 => n21951, C1 => n30486, C2 =>
                           n9486, A => n27376, ZN => n27371);
   U22089 : OAI22_X1 port map( A1 => n25777, A2 => n30480, B1 => n25711, B2 => 
                           n30474, ZN => n27376);
   U22090 : AOI221_X1 port map( B1 => n30492, B2 => n21952, C1 => n30486, C2 =>
                           n9481, A => n27350, ZN => n27345);
   U22091 : OAI22_X1 port map( A1 => n25776, A2 => n30480, B1 => n25710, B2 => 
                           n30474, ZN => n27350);
   U22092 : AOI221_X1 port map( B1 => n30492, B2 => n21953, C1 => n30486, C2 =>
                           n9476, A => n27324, ZN => n27319);
   U22093 : OAI22_X1 port map( A1 => n25775, A2 => n30480, B1 => n25709, B2 => 
                           n30474, ZN => n27324);
   U22094 : AOI221_X1 port map( B1 => n30492, B2 => n21954, C1 => n30486, C2 =>
                           n9471, A => n27298, ZN => n27293);
   U22095 : OAI22_X1 port map( A1 => n25774, A2 => n30480, B1 => n25708, B2 => 
                           n30474, ZN => n27298);
   U22096 : AOI221_X1 port map( B1 => n30492, B2 => n21955, C1 => n30486, C2 =>
                           n9466, A => n27272, ZN => n27267);
   U22097 : OAI22_X1 port map( A1 => n25773, A2 => n30480, B1 => n25707, B2 => 
                           n30474, ZN => n27272);
   U22098 : AOI221_X1 port map( B1 => n30492, B2 => n21956, C1 => n30486, C2 =>
                           n9461, A => n27246, ZN => n27241);
   U22099 : OAI22_X1 port map( A1 => n25772, A2 => n30480, B1 => n25706, B2 => 
                           n30474, ZN => n27246);
   U22100 : AOI221_X1 port map( B1 => n30492, B2 => n21957, C1 => n30486, C2 =>
                           n9456, A => n27220, ZN => n27215);
   U22101 : OAI22_X1 port map( A1 => n25771, A2 => n30480, B1 => n25705, B2 => 
                           n30474, ZN => n27220);
   U22102 : AOI221_X1 port map( B1 => n30492, B2 => n21958, C1 => n30486, C2 =>
                           n9451, A => n27194, ZN => n27189);
   U22103 : OAI22_X1 port map( A1 => n25770, A2 => n30480, B1 => n25704, B2 => 
                           n30474, ZN => n27194);
   U22104 : AOI221_X1 port map( B1 => n30492, B2 => n21959, C1 => n30486, C2 =>
                           n9446, A => n27168, ZN => n27163);
   U22105 : OAI22_X1 port map( A1 => n25769, A2 => n30480, B1 => n25703, B2 => 
                           n30474, ZN => n27168);
   U22106 : AOI221_X1 port map( B1 => n30492, B2 => n21960, C1 => n30486, C2 =>
                           n9441, A => n27142, ZN => n27137);
   U22107 : OAI22_X1 port map( A1 => n25768, A2 => n30480, B1 => n25702, B2 => 
                           n30474, ZN => n27142);
   U22108 : AOI221_X1 port map( B1 => n30492, B2 => n21961, C1 => n30486, C2 =>
                           n9436, A => n27116, ZN => n27111);
   U22109 : OAI22_X1 port map( A1 => n25767, A2 => n30480, B1 => n25701, B2 => 
                           n30474, ZN => n27116);
   U22110 : AOI221_X1 port map( B1 => n30492, B2 => n21962, C1 => n30486, C2 =>
                           n9431, A => n27090, ZN => n27085);
   U22111 : OAI22_X1 port map( A1 => n25766, A2 => n30480, B1 => n25700, B2 => 
                           n30474, ZN => n27090);
   U22112 : AOI221_X1 port map( B1 => n30493, B2 => n21963, C1 => n30487, C2 =>
                           n9426, A => n27064, ZN => n27059);
   U22113 : OAI22_X1 port map( A1 => n25765, A2 => n30481, B1 => n25699, B2 => 
                           n30475, ZN => n27064);
   U22114 : AOI221_X1 port map( B1 => n30493, B2 => n21964, C1 => n30487, C2 =>
                           n9421, A => n27038, ZN => n27033);
   U22115 : OAI22_X1 port map( A1 => n25764, A2 => n30481, B1 => n25698, B2 => 
                           n30475, ZN => n27038);
   U22116 : AOI221_X1 port map( B1 => n30493, B2 => n21965, C1 => n30487, C2 =>
                           n9416, A => n27012, ZN => n27007);
   U22117 : OAI22_X1 port map( A1 => n25763, A2 => n30481, B1 => n25697, B2 => 
                           n30475, ZN => n27012);
   U22118 : AOI221_X1 port map( B1 => n30493, B2 => n21966, C1 => n30487, C2 =>
                           n9411, A => n26986, ZN => n26981);
   U22119 : OAI22_X1 port map( A1 => n25762, A2 => n30481, B1 => n25696, B2 => 
                           n30475, ZN => n26986);
   U22120 : AOI221_X1 port map( B1 => n30493, B2 => n21967, C1 => n30487, C2 =>
                           n9406, A => n26960, ZN => n26955);
   U22121 : OAI22_X1 port map( A1 => n25761, A2 => n30481, B1 => n25695, B2 => 
                           n30475, ZN => n26960);
   U22122 : AOI221_X1 port map( B1 => n30493, B2 => n21968, C1 => n30487, C2 =>
                           n9401, A => n26934, ZN => n26929);
   U22123 : OAI22_X1 port map( A1 => n25760, A2 => n30481, B1 => n25694, B2 => 
                           n30475, ZN => n26934);
   U22124 : AOI221_X1 port map( B1 => n30493, B2 => n21969, C1 => n30487, C2 =>
                           n9396, A => n26908, ZN => n26903);
   U22125 : OAI22_X1 port map( A1 => n25759, A2 => n30481, B1 => n25693, B2 => 
                           n30475, ZN => n26908);
   U22126 : AOI221_X1 port map( B1 => n30493, B2 => n21970, C1 => n30487, C2 =>
                           n9391, A => n26882, ZN => n26877);
   U22127 : OAI22_X1 port map( A1 => n25758, A2 => n30481, B1 => n25692, B2 => 
                           n30475, ZN => n26882);
   U22128 : AOI221_X1 port map( B1 => n30493, B2 => n21971, C1 => n30487, C2 =>
                           n9386, A => n26856, ZN => n26851);
   U22129 : OAI22_X1 port map( A1 => n25757, A2 => n30481, B1 => n25691, B2 => 
                           n30475, ZN => n26856);
   U22130 : AOI221_X1 port map( B1 => n30493, B2 => n21972, C1 => n30487, C2 =>
                           n9381, A => n26830, ZN => n26825);
   U22131 : OAI22_X1 port map( A1 => n25756, A2 => n30481, B1 => n25690, B2 => 
                           n30475, ZN => n26830);
   U22132 : AOI221_X1 port map( B1 => n30493, B2 => n21973, C1 => n30487, C2 =>
                           n9376, A => n26804, ZN => n26799);
   U22133 : OAI22_X1 port map( A1 => n25755, A2 => n30481, B1 => n25689, B2 => 
                           n30475, ZN => n26804);
   U22134 : AOI221_X1 port map( B1 => n30493, B2 => n21974, C1 => n30487, C2 =>
                           n9371, A => n26778, ZN => n26773);
   U22135 : OAI22_X1 port map( A1 => n25754, A2 => n30481, B1 => n25688, B2 => 
                           n30475, ZN => n26778);
   U22136 : AOI221_X1 port map( B1 => n30494, B2 => n21975, C1 => n30488, C2 =>
                           n9366, A => n26752, ZN => n26747);
   U22137 : OAI22_X1 port map( A1 => n25753, A2 => n30482, B1 => n25687, B2 => 
                           n30476, ZN => n26752);
   U22138 : AOI221_X1 port map( B1 => n30494, B2 => n21976, C1 => n30488, C2 =>
                           n9361, A => n26726, ZN => n26721);
   U22139 : OAI22_X1 port map( A1 => n25752, A2 => n30482, B1 => n25686, B2 => 
                           n30476, ZN => n26726);
   U22140 : AOI221_X1 port map( B1 => n30494, B2 => n21977, C1 => n30488, C2 =>
                           n9356, A => n26700, ZN => n26695);
   U22141 : OAI22_X1 port map( A1 => n25751, A2 => n30482, B1 => n25685, B2 => 
                           n30476, ZN => n26700);
   U22142 : AOI221_X1 port map( B1 => n30494, B2 => n21978, C1 => n30488, C2 =>
                           n9351, A => n26674, ZN => n26669);
   U22143 : OAI22_X1 port map( A1 => n25750, A2 => n30482, B1 => n25684, B2 => 
                           n30476, ZN => n26674);
   U22144 : AOI221_X1 port map( B1 => n30494, B2 => n21979, C1 => n30488, C2 =>
                           n9346, A => n26648, ZN => n26643);
   U22145 : OAI22_X1 port map( A1 => n25749, A2 => n30482, B1 => n25683, B2 => 
                           n30476, ZN => n26648);
   U22146 : AOI221_X1 port map( B1 => n30494, B2 => n21980, C1 => n30488, C2 =>
                           n9341, A => n26622, ZN => n26617);
   U22147 : OAI22_X1 port map( A1 => n25748, A2 => n30482, B1 => n25682, B2 => 
                           n30476, ZN => n26622);
   U22148 : AOI221_X1 port map( B1 => n30494, B2 => n21981, C1 => n30488, C2 =>
                           n9336, A => n26596, ZN => n26591);
   U22149 : OAI22_X1 port map( A1 => n25747, A2 => n30482, B1 => n25681, B2 => 
                           n30476, ZN => n26596);
   U22150 : AOI221_X1 port map( B1 => n30494, B2 => n21982, C1 => n30488, C2 =>
                           n9331, A => n26570, ZN => n26565);
   U22151 : OAI22_X1 port map( A1 => n25746, A2 => n30482, B1 => n25680, B2 => 
                           n30476, ZN => n26570);
   U22152 : AOI221_X1 port map( B1 => n30494, B2 => n21983, C1 => n30488, C2 =>
                           n9326, A => n26544, ZN => n26539);
   U22153 : OAI22_X1 port map( A1 => n25745, A2 => n30482, B1 => n25679, B2 => 
                           n30476, ZN => n26544);
   U22154 : AOI221_X1 port map( B1 => n30494, B2 => n21984, C1 => n30488, C2 =>
                           n9321, A => n26518, ZN => n26513);
   U22155 : OAI22_X1 port map( A1 => n25744, A2 => n30482, B1 => n25678, B2 => 
                           n30476, ZN => n26518);
   U22156 : AOI221_X1 port map( B1 => n30494, B2 => n21985, C1 => n30488, C2 =>
                           n9316, A => n26492, ZN => n26487);
   U22157 : OAI22_X1 port map( A1 => n25743, A2 => n30482, B1 => n25677, B2 => 
                           n30476, ZN => n26492);
   U22158 : AOI221_X1 port map( B1 => n30494, B2 => n21986, C1 => n30488, C2 =>
                           n9311, A => n26466, ZN => n26461);
   U22159 : OAI22_X1 port map( A1 => n25742, A2 => n30482, B1 => n25676, B2 => 
                           n30476, ZN => n26466);
   U22160 : AOI221_X1 port map( B1 => n30189, B2 => n29636, C1 => n30183, C2 =>
                           n29444, A => n29304, ZN => n29295);
   U22161 : OAI22_X1 port map( A1 => n9287, A2 => n30177, B1 => n26247, B2 => 
                           n30171, ZN => n29304);
   U22162 : AOI221_X1 port map( B1 => n30189, B2 => n29637, C1 => n30183, C2 =>
                           n29445, A => n29270, ZN => n29265);
   U22163 : OAI22_X1 port map( A1 => n9282, A2 => n30177, B1 => n26246, B2 => 
                           n30171, ZN => n29270);
   U22164 : AOI221_X1 port map( B1 => n30189, B2 => n29638, C1 => n30183, C2 =>
                           n29446, A => n29251, ZN => n29246);
   U22165 : OAI22_X1 port map( A1 => n9277, A2 => n30177, B1 => n26245, B2 => 
                           n30171, ZN => n29251);
   U22166 : AOI221_X1 port map( B1 => n30189, B2 => n29639, C1 => n30183, C2 =>
                           n29447, A => n29232, ZN => n29227);
   U22167 : OAI22_X1 port map( A1 => n9272, A2 => n30177, B1 => n26244, B2 => 
                           n30171, ZN => n29232);
   U22168 : AOI221_X1 port map( B1 => n30189, B2 => n29640, C1 => n30183, C2 =>
                           n29448, A => n29213, ZN => n29208);
   U22169 : OAI22_X1 port map( A1 => n9267, A2 => n30177, B1 => n26243, B2 => 
                           n30171, ZN => n29213);
   U22170 : AOI221_X1 port map( B1 => n30189, B2 => n29641, C1 => n30183, C2 =>
                           n29449, A => n29194, ZN => n29189);
   U22171 : OAI22_X1 port map( A1 => n9262, A2 => n30177, B1 => n26242, B2 => 
                           n30171, ZN => n29194);
   U22172 : AOI221_X1 port map( B1 => n30189, B2 => n29642, C1 => n30183, C2 =>
                           n29450, A => n29175, ZN => n29170);
   U22173 : OAI22_X1 port map( A1 => n9257, A2 => n30177, B1 => n26241, B2 => 
                           n30171, ZN => n29175);
   U22174 : AOI221_X1 port map( B1 => n30189, B2 => n29643, C1 => n30183, C2 =>
                           n29451, A => n29156, ZN => n29151);
   U22175 : OAI22_X1 port map( A1 => n9252, A2 => n30177, B1 => n26240, B2 => 
                           n30171, ZN => n29156);
   U22176 : AOI221_X1 port map( B1 => n30189, B2 => n29644, C1 => n30183, C2 =>
                           n29452, A => n29137, ZN => n29132);
   U22177 : OAI22_X1 port map( A1 => n9247, A2 => n30177, B1 => n26239, B2 => 
                           n30171, ZN => n29137);
   U22178 : AOI221_X1 port map( B1 => n30189, B2 => n29645, C1 => n30183, C2 =>
                           n29453, A => n29118, ZN => n29113);
   U22179 : OAI22_X1 port map( A1 => n9242, A2 => n30177, B1 => n26238, B2 => 
                           n30171, ZN => n29118);
   U22180 : AOI221_X1 port map( B1 => n30189, B2 => n29646, C1 => n30183, C2 =>
                           n29454, A => n29099, ZN => n29094);
   U22181 : OAI22_X1 port map( A1 => n9237, A2 => n30177, B1 => n26237, B2 => 
                           n30171, ZN => n29099);
   U22182 : AOI221_X1 port map( B1 => n30189, B2 => n29647, C1 => n30183, C2 =>
                           n29455, A => n29080, ZN => n29075);
   U22183 : OAI22_X1 port map( A1 => n9232, A2 => n30177, B1 => n26236, B2 => 
                           n30171, ZN => n29080);
   U22184 : AOI221_X1 port map( B1 => n30190, B2 => n29648, C1 => n30184, C2 =>
                           n29456, A => n29061, ZN => n29056);
   U22185 : OAI22_X1 port map( A1 => n9227, A2 => n30178, B1 => n9995, B2 => 
                           n30172, ZN => n29061);
   U22186 : AOI221_X1 port map( B1 => n30190, B2 => n29649, C1 => n30184, C2 =>
                           n29457, A => n29042, ZN => n29037);
   U22187 : OAI22_X1 port map( A1 => n9222, A2 => n30178, B1 => n9990, B2 => 
                           n30172, ZN => n29042);
   U22188 : AOI221_X1 port map( B1 => n30190, B2 => n29650, C1 => n30184, C2 =>
                           n29458, A => n29023, ZN => n29018);
   U22189 : OAI22_X1 port map( A1 => n9217, A2 => n30178, B1 => n9985, B2 => 
                           n30172, ZN => n29023);
   U22190 : AOI221_X1 port map( B1 => n30190, B2 => n29651, C1 => n30184, C2 =>
                           n29459, A => n29004, ZN => n28999);
   U22191 : OAI22_X1 port map( A1 => n9212, A2 => n30178, B1 => n9980, B2 => 
                           n30172, ZN => n29004);
   U22192 : AOI221_X1 port map( B1 => n30190, B2 => n29652, C1 => n30184, C2 =>
                           n29460, A => n28985, ZN => n28980);
   U22193 : OAI22_X1 port map( A1 => n9207, A2 => n30178, B1 => n9975, B2 => 
                           n30172, ZN => n28985);
   U22194 : AOI221_X1 port map( B1 => n30190, B2 => n29653, C1 => n30184, C2 =>
                           n29461, A => n28966, ZN => n28961);
   U22195 : OAI22_X1 port map( A1 => n9202, A2 => n30178, B1 => n9970, B2 => 
                           n30172, ZN => n28966);
   U22196 : AOI221_X1 port map( B1 => n30190, B2 => n29654, C1 => n30184, C2 =>
                           n29462, A => n28947, ZN => n28942);
   U22197 : OAI22_X1 port map( A1 => n9197, A2 => n30178, B1 => n9965, B2 => 
                           n30172, ZN => n28947);
   U22198 : AOI221_X1 port map( B1 => n30190, B2 => n29655, C1 => n30184, C2 =>
                           n29463, A => n28928, ZN => n28923);
   U22199 : OAI22_X1 port map( A1 => n9192, A2 => n30178, B1 => n9960, B2 => 
                           n30172, ZN => n28928);
   U22200 : AOI221_X1 port map( B1 => n30190, B2 => n29656, C1 => n30184, C2 =>
                           n29464, A => n28909, ZN => n28904);
   U22201 : OAI22_X1 port map( A1 => n9187, A2 => n30178, B1 => n9955, B2 => 
                           n30172, ZN => n28909);
   U22202 : AOI221_X1 port map( B1 => n30190, B2 => n29657, C1 => n30184, C2 =>
                           n29465, A => n28890, ZN => n28885);
   U22203 : OAI22_X1 port map( A1 => n9182, A2 => n30178, B1 => n9950, B2 => 
                           n30172, ZN => n28890);
   U22204 : AOI221_X1 port map( B1 => n30190, B2 => n29658, C1 => n30184, C2 =>
                           n29466, A => n28871, ZN => n28866);
   U22205 : OAI22_X1 port map( A1 => n9177, A2 => n30178, B1 => n9945, B2 => 
                           n30172, ZN => n28871);
   U22206 : AOI221_X1 port map( B1 => n30190, B2 => n29659, C1 => n30184, C2 =>
                           n29467, A => n28852, ZN => n28847);
   U22207 : OAI22_X1 port map( A1 => n9172, A2 => n30178, B1 => n9940, B2 => 
                           n30172, ZN => n28852);
   U22208 : AOI221_X1 port map( B1 => n30191, B2 => n29660, C1 => n30185, C2 =>
                           n29468, A => n28833, ZN => n28828);
   U22209 : OAI22_X1 port map( A1 => n9167, A2 => n30179, B1 => n9935, B2 => 
                           n30173, ZN => n28833);
   U22210 : AOI221_X1 port map( B1 => n30191, B2 => n29661, C1 => n30185, C2 =>
                           n29469, A => n28814, ZN => n28809);
   U22211 : OAI22_X1 port map( A1 => n9162, A2 => n30179, B1 => n9930, B2 => 
                           n30173, ZN => n28814);
   U22212 : AOI221_X1 port map( B1 => n30191, B2 => n29662, C1 => n30185, C2 =>
                           n29470, A => n28795, ZN => n28790);
   U22213 : OAI22_X1 port map( A1 => n9157, A2 => n30179, B1 => n9925, B2 => 
                           n30173, ZN => n28795);
   U22214 : AOI221_X1 port map( B1 => n30191, B2 => n29663, C1 => n30185, C2 =>
                           n29471, A => n28776, ZN => n28771);
   U22215 : OAI22_X1 port map( A1 => n9152, A2 => n30179, B1 => n9920, B2 => 
                           n30173, ZN => n28776);
   U22216 : AOI221_X1 port map( B1 => n30191, B2 => n29664, C1 => n30185, C2 =>
                           n29472, A => n28757, ZN => n28752);
   U22217 : OAI22_X1 port map( A1 => n9147, A2 => n30179, B1 => n9915, B2 => 
                           n30173, ZN => n28757);
   U22218 : AOI221_X1 port map( B1 => n30191, B2 => n29665, C1 => n30185, C2 =>
                           n29473, A => n28738, ZN => n28733);
   U22219 : OAI22_X1 port map( A1 => n9142, A2 => n30179, B1 => n9910, B2 => 
                           n30173, ZN => n28738);
   U22220 : AOI221_X1 port map( B1 => n30191, B2 => n29666, C1 => n30185, C2 =>
                           n29474, A => n28719, ZN => n28714);
   U22221 : OAI22_X1 port map( A1 => n9137, A2 => n30179, B1 => n9905, B2 => 
                           n30173, ZN => n28719);
   U22222 : AOI221_X1 port map( B1 => n30191, B2 => n29667, C1 => n30185, C2 =>
                           n29475, A => n28700, ZN => n28695);
   U22223 : OAI22_X1 port map( A1 => n9132, A2 => n30179, B1 => n9900, B2 => 
                           n30173, ZN => n28700);
   U22224 : AOI221_X1 port map( B1 => n30191, B2 => n29668, C1 => n30185, C2 =>
                           n29476, A => n28681, ZN => n28676);
   U22225 : OAI22_X1 port map( A1 => n9127, A2 => n30179, B1 => n9895, B2 => 
                           n30173, ZN => n28681);
   U22226 : AOI221_X1 port map( B1 => n30191, B2 => n29669, C1 => n30185, C2 =>
                           n29477, A => n28662, ZN => n28657);
   U22227 : OAI22_X1 port map( A1 => n9122, A2 => n30179, B1 => n9890, B2 => 
                           n30173, ZN => n28662);
   U22228 : AOI221_X1 port map( B1 => n30191, B2 => n29670, C1 => n30185, C2 =>
                           n29478, A => n28643, ZN => n28638);
   U22229 : OAI22_X1 port map( A1 => n9117, A2 => n30179, B1 => n9885, B2 => 
                           n30173, ZN => n28643);
   U22230 : AOI221_X1 port map( B1 => n30191, B2 => n29671, C1 => n30185, C2 =>
                           n29479, A => n28624, ZN => n28619);
   U22231 : OAI22_X1 port map( A1 => n9112, A2 => n30179, B1 => n9880, B2 => 
                           n30173, ZN => n28624);
   U22232 : AOI221_X1 port map( B1 => n30192, B2 => n29672, C1 => n30186, C2 =>
                           n29480, A => n28605, ZN => n28600);
   U22233 : OAI22_X1 port map( A1 => n9107, A2 => n30180, B1 => n9875, B2 => 
                           n30174, ZN => n28605);
   U22234 : AOI221_X1 port map( B1 => n30192, B2 => n29673, C1 => n30186, C2 =>
                           n29481, A => n28586, ZN => n28581);
   U22235 : OAI22_X1 port map( A1 => n9102, A2 => n30180, B1 => n9870, B2 => 
                           n30174, ZN => n28586);
   U22236 : AOI221_X1 port map( B1 => n30192, B2 => n29674, C1 => n30186, C2 =>
                           n29482, A => n28567, ZN => n28562);
   U22237 : OAI22_X1 port map( A1 => n9097, A2 => n30180, B1 => n9865, B2 => 
                           n30174, ZN => n28567);
   U22238 : AOI221_X1 port map( B1 => n30192, B2 => n29675, C1 => n30186, C2 =>
                           n29483, A => n28548, ZN => n28543);
   U22239 : OAI22_X1 port map( A1 => n9092, A2 => n30180, B1 => n9860, B2 => 
                           n30174, ZN => n28548);
   U22240 : AOI221_X1 port map( B1 => n30192, B2 => n29676, C1 => n30186, C2 =>
                           n29484, A => n28529, ZN => n28524);
   U22241 : OAI22_X1 port map( A1 => n9087, A2 => n30180, B1 => n9855, B2 => 
                           n30174, ZN => n28529);
   U22242 : AOI221_X1 port map( B1 => n30192, B2 => n29677, C1 => n30186, C2 =>
                           n29485, A => n28510, ZN => n28505);
   U22243 : OAI22_X1 port map( A1 => n9082, A2 => n30180, B1 => n9850, B2 => 
                           n30174, ZN => n28510);
   U22244 : AOI221_X1 port map( B1 => n30192, B2 => n29678, C1 => n30186, C2 =>
                           n29486, A => n28491, ZN => n28486);
   U22245 : OAI22_X1 port map( A1 => n9077, A2 => n30180, B1 => n9845, B2 => 
                           n30174, ZN => n28491);
   U22246 : AOI221_X1 port map( B1 => n30192, B2 => n29679, C1 => n30186, C2 =>
                           n29487, A => n28472, ZN => n28467);
   U22247 : OAI22_X1 port map( A1 => n9072, A2 => n30180, B1 => n9840, B2 => 
                           n30174, ZN => n28472);
   U22248 : AOI221_X1 port map( B1 => n30192, B2 => n29680, C1 => n30186, C2 =>
                           n29488, A => n28453, ZN => n28448);
   U22249 : OAI22_X1 port map( A1 => n9067, A2 => n30180, B1 => n9835, B2 => 
                           n30174, ZN => n28453);
   U22250 : AOI221_X1 port map( B1 => n30192, B2 => n29681, C1 => n30186, C2 =>
                           n29489, A => n28434, ZN => n28429);
   U22251 : OAI22_X1 port map( A1 => n9062, A2 => n30180, B1 => n9830, B2 => 
                           n30174, ZN => n28434);
   U22252 : AOI221_X1 port map( B1 => n30192, B2 => n29682, C1 => n30186, C2 =>
                           n29490, A => n28415, ZN => n28410);
   U22253 : OAI22_X1 port map( A1 => n9057, A2 => n30180, B1 => n9825, B2 => 
                           n30174, ZN => n28415);
   U22254 : AOI221_X1 port map( B1 => n30192, B2 => n29683, C1 => n30186, C2 =>
                           n29491, A => n28396, ZN => n28391);
   U22255 : OAI22_X1 port map( A1 => n9052, A2 => n30180, B1 => n9820, B2 => 
                           n30174, ZN => n28396);
   U22256 : AOI221_X1 port map( B1 => n30193, B2 => n29684, C1 => n30187, C2 =>
                           n29492, A => n28377, ZN => n28372);
   U22257 : OAI22_X1 port map( A1 => n9047, A2 => n30181, B1 => n9815, B2 => 
                           n30175, ZN => n28377);
   U22258 : AOI221_X1 port map( B1 => n30193, B2 => n29685, C1 => n30187, C2 =>
                           n29493, A => n28358, ZN => n28353);
   U22259 : OAI22_X1 port map( A1 => n9042, A2 => n30181, B1 => n9810, B2 => 
                           n30175, ZN => n28358);
   U22260 : AOI221_X1 port map( B1 => n30193, B2 => n29686, C1 => n30187, C2 =>
                           n29494, A => n28339, ZN => n28334);
   U22261 : OAI22_X1 port map( A1 => n9037, A2 => n30181, B1 => n9805, B2 => 
                           n30175, ZN => n28339);
   U22262 : AOI221_X1 port map( B1 => n30193, B2 => n29687, C1 => n30187, C2 =>
                           n29495, A => n28320, ZN => n28315);
   U22263 : OAI22_X1 port map( A1 => n9032, A2 => n30181, B1 => n9800, B2 => 
                           n30175, ZN => n28320);
   U22264 : AOI221_X1 port map( B1 => n30193, B2 => n29688, C1 => n30187, C2 =>
                           n29496, A => n28301, ZN => n28296);
   U22265 : OAI22_X1 port map( A1 => n9027, A2 => n30181, B1 => n9795, B2 => 
                           n30175, ZN => n28301);
   U22266 : AOI221_X1 port map( B1 => n30193, B2 => n29689, C1 => n30187, C2 =>
                           n29497, A => n28282, ZN => n28277);
   U22267 : OAI22_X1 port map( A1 => n9022, A2 => n30181, B1 => n9790, B2 => 
                           n30175, ZN => n28282);
   U22268 : AOI221_X1 port map( B1 => n30193, B2 => n29690, C1 => n30187, C2 =>
                           n29498, A => n28263, ZN => n28258);
   U22269 : OAI22_X1 port map( A1 => n9017, A2 => n30181, B1 => n9785, B2 => 
                           n30175, ZN => n28263);
   U22270 : AOI221_X1 port map( B1 => n30193, B2 => n29691, C1 => n30187, C2 =>
                           n29499, A => n28244, ZN => n28239);
   U22271 : OAI22_X1 port map( A1 => n9012, A2 => n30181, B1 => n9780, B2 => 
                           n30175, ZN => n28244);
   U22272 : AOI221_X1 port map( B1 => n30193, B2 => n29692, C1 => n30187, C2 =>
                           n29500, A => n28225, ZN => n28220);
   U22273 : OAI22_X1 port map( A1 => n9007, A2 => n30181, B1 => n9775, B2 => 
                           n30175, ZN => n28225);
   U22274 : AOI221_X1 port map( B1 => n30193, B2 => n29693, C1 => n30187, C2 =>
                           n29501, A => n28206, ZN => n28201);
   U22275 : OAI22_X1 port map( A1 => n9002, A2 => n30181, B1 => n9770, B2 => 
                           n30175, ZN => n28206);
   U22276 : AOI221_X1 port map( B1 => n30193, B2 => n29694, C1 => n30187, C2 =>
                           n29502, A => n28187, ZN => n28182);
   U22277 : OAI22_X1 port map( A1 => n8997, A2 => n30181, B1 => n9765, B2 => 
                           n30175, ZN => n28187);
   U22278 : AOI221_X1 port map( B1 => n30193, B2 => n29695, C1 => n30187, C2 =>
                           n29503, A => n28168, ZN => n28163);
   U22279 : OAI22_X1 port map( A1 => n8992, A2 => n30181, B1 => n9760, B2 => 
                           n30175, ZN => n28168);
   U22280 : AOI221_X1 port map( B1 => n30194, B2 => n29696, C1 => n30188, C2 =>
                           n29504, A => n28149, ZN => n28144);
   U22281 : OAI22_X1 port map( A1 => n8987, A2 => n30182, B1 => n9755, B2 => 
                           n30176, ZN => n28149);
   U22282 : AOI221_X1 port map( B1 => n30290, B2 => n22239, C1 => n30284, C2 =>
                           n9676, A => n28141, ZN => n28136);
   U22283 : OAI22_X1 port map( A1 => n9612, A2 => n30278, B1 => n17776, B2 => 
                           n30272, ZN => n28141);
   U22284 : AOI221_X1 port map( B1 => n30194, B2 => n29697, C1 => n30188, C2 =>
                           n29505, A => n28130, ZN => n28125);
   U22285 : OAI22_X1 port map( A1 => n8982, A2 => n30182, B1 => n9750, B2 => 
                           n30176, ZN => n28130);
   U22286 : AOI221_X1 port map( B1 => n30290, B2 => n22240, C1 => n30284, C2 =>
                           n9675, A => n28122, ZN => n28117);
   U22287 : OAI22_X1 port map( A1 => n9611, A2 => n30278, B1 => n17775, B2 => 
                           n30272, ZN => n28122);
   U22288 : AOI221_X1 port map( B1 => n30194, B2 => n29698, C1 => n30188, C2 =>
                           n29506, A => n28111, ZN => n28106);
   U22289 : OAI22_X1 port map( A1 => n8977, A2 => n30182, B1 => n9745, B2 => 
                           n30176, ZN => n28111);
   U22290 : AOI221_X1 port map( B1 => n30290, B2 => n22241, C1 => n30284, C2 =>
                           n9674, A => n28103, ZN => n28098);
   U22291 : OAI22_X1 port map( A1 => n9610, A2 => n30278, B1 => n17774, B2 => 
                           n30272, ZN => n28103);
   U22292 : AOI221_X1 port map( B1 => n30194, B2 => n29699, C1 => n30188, C2 =>
                           n29507, A => n28085, ZN => n28070);
   U22293 : OAI22_X1 port map( A1 => n8972, A2 => n30182, B1 => n9740, B2 => 
                           n30176, ZN => n28085);
   U22294 : AOI221_X1 port map( B1 => n30290, B2 => n22242, C1 => n30284, C2 =>
                           n9673, A => n28061, ZN => n28046);
   U22295 : OAI22_X1 port map( A1 => n9609, A2 => n30278, B1 => n17772, B2 => 
                           n30272, ZN => n28061);
   U22296 : AOI221_X1 port map( B1 => n30393, B2 => n29636, C1 => n30387, C2 =>
                           n29444, A => n28027, ZN => n28015);
   U22297 : OAI22_X1 port map( A1 => n9287, A2 => n30381, B1 => n26247, B2 => 
                           n30375, ZN => n28027);
   U22298 : AOI221_X1 port map( B1 => n30393, B2 => n29637, C1 => n30387, C2 =>
                           n29445, A => n27986, ZN => n27977);
   U22299 : OAI22_X1 port map( A1 => n9282, A2 => n30381, B1 => n26246, B2 => 
                           n30375, ZN => n27986);
   U22300 : AOI221_X1 port map( B1 => n30393, B2 => n29638, C1 => n30387, C2 =>
                           n29446, A => n27960, ZN => n27951);
   U22301 : OAI22_X1 port map( A1 => n9277, A2 => n30381, B1 => n26245, B2 => 
                           n30375, ZN => n27960);
   U22302 : AOI221_X1 port map( B1 => n30393, B2 => n29639, C1 => n30387, C2 =>
                           n29447, A => n27934, ZN => n27925);
   U22303 : OAI22_X1 port map( A1 => n9272, A2 => n30381, B1 => n26244, B2 => 
                           n30375, ZN => n27934);
   U22304 : AOI221_X1 port map( B1 => n30393, B2 => n29640, C1 => n30387, C2 =>
                           n29448, A => n27908, ZN => n27899);
   U22305 : OAI22_X1 port map( A1 => n9267, A2 => n30381, B1 => n26243, B2 => 
                           n30375, ZN => n27908);
   U22306 : AOI221_X1 port map( B1 => n30393, B2 => n29641, C1 => n30387, C2 =>
                           n29449, A => n27882, ZN => n27873);
   U22307 : OAI22_X1 port map( A1 => n9262, A2 => n30381, B1 => n26242, B2 => 
                           n30375, ZN => n27882);
   U22308 : AOI221_X1 port map( B1 => n30393, B2 => n29642, C1 => n30387, C2 =>
                           n29450, A => n27856, ZN => n27847);
   U22309 : OAI22_X1 port map( A1 => n9257, A2 => n30381, B1 => n26241, B2 => 
                           n30375, ZN => n27856);
   U22310 : AOI221_X1 port map( B1 => n30393, B2 => n29643, C1 => n30387, C2 =>
                           n29451, A => n27830, ZN => n27821);
   U22311 : OAI22_X1 port map( A1 => n9252, A2 => n30381, B1 => n26240, B2 => 
                           n30375, ZN => n27830);
   U22312 : AOI221_X1 port map( B1 => n30393, B2 => n29644, C1 => n30387, C2 =>
                           n29452, A => n27804, ZN => n27795);
   U22313 : OAI22_X1 port map( A1 => n9247, A2 => n30381, B1 => n26239, B2 => 
                           n30375, ZN => n27804);
   U22314 : AOI221_X1 port map( B1 => n30393, B2 => n29645, C1 => n30387, C2 =>
                           n29453, A => n27778, ZN => n27769);
   U22315 : OAI22_X1 port map( A1 => n9242, A2 => n30381, B1 => n26238, B2 => 
                           n30375, ZN => n27778);
   U22316 : AOI221_X1 port map( B1 => n30393, B2 => n29646, C1 => n30387, C2 =>
                           n29454, A => n27752, ZN => n27743);
   U22317 : OAI22_X1 port map( A1 => n9237, A2 => n30381, B1 => n26237, B2 => 
                           n30375, ZN => n27752);
   U22318 : AOI221_X1 port map( B1 => n30393, B2 => n29647, C1 => n30387, C2 =>
                           n29455, A => n27726, ZN => n27717);
   U22319 : OAI22_X1 port map( A1 => n9232, A2 => n30381, B1 => n26236, B2 => 
                           n30375, ZN => n27726);
   U22320 : AOI221_X1 port map( B1 => n30394, B2 => n29648, C1 => n30388, C2 =>
                           n29456, A => n27700, ZN => n27691);
   U22321 : OAI22_X1 port map( A1 => n9227, A2 => n30382, B1 => n9995, B2 => 
                           n30376, ZN => n27700);
   U22322 : AOI221_X1 port map( B1 => n30394, B2 => n29649, C1 => n30388, C2 =>
                           n29457, A => n27674, ZN => n27665);
   U22323 : OAI22_X1 port map( A1 => n9222, A2 => n30382, B1 => n9990, B2 => 
                           n30376, ZN => n27674);
   U22324 : AOI221_X1 port map( B1 => n30394, B2 => n29650, C1 => n30388, C2 =>
                           n29458, A => n27648, ZN => n27639);
   U22325 : OAI22_X1 port map( A1 => n9217, A2 => n30382, B1 => n9985, B2 => 
                           n30376, ZN => n27648);
   U22326 : AOI221_X1 port map( B1 => n30394, B2 => n29651, C1 => n30388, C2 =>
                           n29459, A => n27622, ZN => n27613);
   U22327 : OAI22_X1 port map( A1 => n9212, A2 => n30382, B1 => n9980, B2 => 
                           n30376, ZN => n27622);
   U22328 : AOI221_X1 port map( B1 => n30394, B2 => n29652, C1 => n30388, C2 =>
                           n29460, A => n27596, ZN => n27587);
   U22329 : OAI22_X1 port map( A1 => n9207, A2 => n30382, B1 => n9975, B2 => 
                           n30376, ZN => n27596);
   U22330 : AOI221_X1 port map( B1 => n30394, B2 => n29653, C1 => n30388, C2 =>
                           n29461, A => n27570, ZN => n27561);
   U22331 : OAI22_X1 port map( A1 => n9202, A2 => n30382, B1 => n9970, B2 => 
                           n30376, ZN => n27570);
   U22332 : AOI221_X1 port map( B1 => n30394, B2 => n29654, C1 => n30388, C2 =>
                           n29462, A => n27544, ZN => n27535);
   U22333 : OAI22_X1 port map( A1 => n9197, A2 => n30382, B1 => n9965, B2 => 
                           n30376, ZN => n27544);
   U22334 : AOI221_X1 port map( B1 => n30394, B2 => n29655, C1 => n30388, C2 =>
                           n29463, A => n27518, ZN => n27509);
   U22335 : OAI22_X1 port map( A1 => n9192, A2 => n30382, B1 => n9960, B2 => 
                           n30376, ZN => n27518);
   U22336 : AOI221_X1 port map( B1 => n30394, B2 => n29656, C1 => n30388, C2 =>
                           n29464, A => n27492, ZN => n27483);
   U22337 : OAI22_X1 port map( A1 => n9187, A2 => n30382, B1 => n9955, B2 => 
                           n30376, ZN => n27492);
   U22338 : AOI221_X1 port map( B1 => n30394, B2 => n29657, C1 => n30388, C2 =>
                           n29465, A => n27466, ZN => n27457);
   U22339 : OAI22_X1 port map( A1 => n9182, A2 => n30382, B1 => n9950, B2 => 
                           n30376, ZN => n27466);
   U22340 : AOI221_X1 port map( B1 => n30394, B2 => n29658, C1 => n30388, C2 =>
                           n29466, A => n27440, ZN => n27431);
   U22341 : OAI22_X1 port map( A1 => n9177, A2 => n30382, B1 => n9945, B2 => 
                           n30376, ZN => n27440);
   U22342 : AOI221_X1 port map( B1 => n30394, B2 => n29659, C1 => n30388, C2 =>
                           n29467, A => n27414, ZN => n27405);
   U22343 : OAI22_X1 port map( A1 => n9172, A2 => n30382, B1 => n9940, B2 => 
                           n30376, ZN => n27414);
   U22344 : AOI221_X1 port map( B1 => n30395, B2 => n29660, C1 => n30389, C2 =>
                           n29468, A => n27388, ZN => n27379);
   U22345 : OAI22_X1 port map( A1 => n9167, A2 => n30383, B1 => n9935, B2 => 
                           n30377, ZN => n27388);
   U22346 : AOI221_X1 port map( B1 => n30395, B2 => n29661, C1 => n30389, C2 =>
                           n29469, A => n27362, ZN => n27353);
   U22347 : OAI22_X1 port map( A1 => n9162, A2 => n30383, B1 => n9930, B2 => 
                           n30377, ZN => n27362);
   U22348 : AOI221_X1 port map( B1 => n30395, B2 => n29662, C1 => n30389, C2 =>
                           n29470, A => n27336, ZN => n27327);
   U22349 : OAI22_X1 port map( A1 => n9157, A2 => n30383, B1 => n9925, B2 => 
                           n30377, ZN => n27336);
   U22350 : AOI221_X1 port map( B1 => n30395, B2 => n29663, C1 => n30389, C2 =>
                           n29471, A => n27310, ZN => n27301);
   U22351 : OAI22_X1 port map( A1 => n9152, A2 => n30383, B1 => n9920, B2 => 
                           n30377, ZN => n27310);
   U22352 : AOI221_X1 port map( B1 => n30395, B2 => n29664, C1 => n30389, C2 =>
                           n29472, A => n27284, ZN => n27275);
   U22353 : OAI22_X1 port map( A1 => n9147, A2 => n30383, B1 => n9915, B2 => 
                           n30377, ZN => n27284);
   U22354 : AOI221_X1 port map( B1 => n30395, B2 => n29665, C1 => n30389, C2 =>
                           n29473, A => n27258, ZN => n27249);
   U22355 : OAI22_X1 port map( A1 => n9142, A2 => n30383, B1 => n9910, B2 => 
                           n30377, ZN => n27258);
   U22356 : AOI221_X1 port map( B1 => n30395, B2 => n29666, C1 => n30389, C2 =>
                           n29474, A => n27232, ZN => n27223);
   U22357 : OAI22_X1 port map( A1 => n9137, A2 => n30383, B1 => n9905, B2 => 
                           n30377, ZN => n27232);
   U22358 : AOI221_X1 port map( B1 => n30395, B2 => n29667, C1 => n30389, C2 =>
                           n29475, A => n27206, ZN => n27197);
   U22359 : OAI22_X1 port map( A1 => n9132, A2 => n30383, B1 => n9900, B2 => 
                           n30377, ZN => n27206);
   U22360 : AOI221_X1 port map( B1 => n30395, B2 => n29668, C1 => n30389, C2 =>
                           n29476, A => n27180, ZN => n27171);
   U22361 : OAI22_X1 port map( A1 => n9127, A2 => n30383, B1 => n9895, B2 => 
                           n30377, ZN => n27180);
   U22362 : AOI221_X1 port map( B1 => n30395, B2 => n29669, C1 => n30389, C2 =>
                           n29477, A => n27154, ZN => n27145);
   U22363 : OAI22_X1 port map( A1 => n9122, A2 => n30383, B1 => n9890, B2 => 
                           n30377, ZN => n27154);
   U22364 : AOI221_X1 port map( B1 => n30395, B2 => n29670, C1 => n30389, C2 =>
                           n29478, A => n27128, ZN => n27119);
   U22365 : OAI22_X1 port map( A1 => n9117, A2 => n30383, B1 => n9885, B2 => 
                           n30377, ZN => n27128);
   U22366 : AOI221_X1 port map( B1 => n30395, B2 => n29671, C1 => n30389, C2 =>
                           n29479, A => n27102, ZN => n27093);
   U22367 : OAI22_X1 port map( A1 => n9112, A2 => n30383, B1 => n9880, B2 => 
                           n30377, ZN => n27102);
   U22368 : AOI221_X1 port map( B1 => n30396, B2 => n29672, C1 => n30390, C2 =>
                           n29480, A => n27076, ZN => n27067);
   U22369 : OAI22_X1 port map( A1 => n9107, A2 => n30384, B1 => n9875, B2 => 
                           n30378, ZN => n27076);
   U22370 : AOI221_X1 port map( B1 => n30396, B2 => n29673, C1 => n30390, C2 =>
                           n29481, A => n27050, ZN => n27041);
   U22371 : OAI22_X1 port map( A1 => n9102, A2 => n30384, B1 => n9870, B2 => 
                           n30378, ZN => n27050);
   U22372 : AOI221_X1 port map( B1 => n30396, B2 => n29674, C1 => n30390, C2 =>
                           n29482, A => n27024, ZN => n27015);
   U22373 : OAI22_X1 port map( A1 => n9097, A2 => n30384, B1 => n9865, B2 => 
                           n30378, ZN => n27024);
   U22374 : AOI221_X1 port map( B1 => n30396, B2 => n29675, C1 => n30390, C2 =>
                           n29483, A => n26998, ZN => n26989);
   U22375 : OAI22_X1 port map( A1 => n9092, A2 => n30384, B1 => n9860, B2 => 
                           n30378, ZN => n26998);
   U22376 : AOI221_X1 port map( B1 => n30396, B2 => n29676, C1 => n30390, C2 =>
                           n29484, A => n26972, ZN => n26963);
   U22377 : OAI22_X1 port map( A1 => n9087, A2 => n30384, B1 => n9855, B2 => 
                           n30378, ZN => n26972);
   U22378 : AOI221_X1 port map( B1 => n30396, B2 => n29677, C1 => n30390, C2 =>
                           n29485, A => n26946, ZN => n26937);
   U22379 : OAI22_X1 port map( A1 => n9082, A2 => n30384, B1 => n9850, B2 => 
                           n30378, ZN => n26946);
   U22380 : AOI221_X1 port map( B1 => n30396, B2 => n29678, C1 => n30390, C2 =>
                           n29486, A => n26920, ZN => n26911);
   U22381 : OAI22_X1 port map( A1 => n9077, A2 => n30384, B1 => n9845, B2 => 
                           n30378, ZN => n26920);
   U22382 : AOI221_X1 port map( B1 => n30396, B2 => n29679, C1 => n30390, C2 =>
                           n29487, A => n26894, ZN => n26885);
   U22383 : OAI22_X1 port map( A1 => n9072, A2 => n30384, B1 => n9840, B2 => 
                           n30378, ZN => n26894);
   U22384 : AOI221_X1 port map( B1 => n30396, B2 => n29680, C1 => n30390, C2 =>
                           n29488, A => n26868, ZN => n26859);
   U22385 : OAI22_X1 port map( A1 => n9067, A2 => n30384, B1 => n9835, B2 => 
                           n30378, ZN => n26868);
   U22386 : AOI221_X1 port map( B1 => n30396, B2 => n29681, C1 => n30390, C2 =>
                           n29489, A => n26842, ZN => n26833);
   U22387 : OAI22_X1 port map( A1 => n9062, A2 => n30384, B1 => n9830, B2 => 
                           n30378, ZN => n26842);
   U22388 : AOI221_X1 port map( B1 => n30396, B2 => n29682, C1 => n30390, C2 =>
                           n29490, A => n26816, ZN => n26807);
   U22389 : OAI22_X1 port map( A1 => n9057, A2 => n30384, B1 => n9825, B2 => 
                           n30378, ZN => n26816);
   U22390 : AOI221_X1 port map( B1 => n30396, B2 => n29683, C1 => n30390, C2 =>
                           n29491, A => n26790, ZN => n26781);
   U22391 : OAI22_X1 port map( A1 => n9052, A2 => n30384, B1 => n9820, B2 => 
                           n30378, ZN => n26790);
   U22392 : AOI221_X1 port map( B1 => n30397, B2 => n29684, C1 => n30391, C2 =>
                           n29492, A => n26764, ZN => n26755);
   U22393 : OAI22_X1 port map( A1 => n9047, A2 => n30385, B1 => n9815, B2 => 
                           n30379, ZN => n26764);
   U22394 : AOI221_X1 port map( B1 => n30397, B2 => n29685, C1 => n30391, C2 =>
                           n29493, A => n26738, ZN => n26729);
   U22395 : OAI22_X1 port map( A1 => n9042, A2 => n30385, B1 => n9810, B2 => 
                           n30379, ZN => n26738);
   U22396 : AOI221_X1 port map( B1 => n30397, B2 => n29686, C1 => n30391, C2 =>
                           n29494, A => n26712, ZN => n26703);
   U22397 : OAI22_X1 port map( A1 => n9037, A2 => n30385, B1 => n9805, B2 => 
                           n30379, ZN => n26712);
   U22398 : AOI221_X1 port map( B1 => n30397, B2 => n29687, C1 => n30391, C2 =>
                           n29495, A => n26686, ZN => n26677);
   U22399 : OAI22_X1 port map( A1 => n9032, A2 => n30385, B1 => n9800, B2 => 
                           n30379, ZN => n26686);
   U22400 : AOI221_X1 port map( B1 => n30397, B2 => n29688, C1 => n30391, C2 =>
                           n29496, A => n26660, ZN => n26651);
   U22401 : OAI22_X1 port map( A1 => n9027, A2 => n30385, B1 => n9795, B2 => 
                           n30379, ZN => n26660);
   U22402 : AOI221_X1 port map( B1 => n30397, B2 => n29689, C1 => n30391, C2 =>
                           n29497, A => n26634, ZN => n26625);
   U22403 : OAI22_X1 port map( A1 => n9022, A2 => n30385, B1 => n9790, B2 => 
                           n30379, ZN => n26634);
   U22404 : AOI221_X1 port map( B1 => n30397, B2 => n29690, C1 => n30391, C2 =>
                           n29498, A => n26608, ZN => n26599);
   U22405 : OAI22_X1 port map( A1 => n9017, A2 => n30385, B1 => n9785, B2 => 
                           n30379, ZN => n26608);
   U22406 : AOI221_X1 port map( B1 => n30397, B2 => n29691, C1 => n30391, C2 =>
                           n29499, A => n26582, ZN => n26573);
   U22407 : OAI22_X1 port map( A1 => n9012, A2 => n30385, B1 => n9780, B2 => 
                           n30379, ZN => n26582);
   U22408 : AOI221_X1 port map( B1 => n30397, B2 => n29692, C1 => n30391, C2 =>
                           n29500, A => n26556, ZN => n26547);
   U22409 : OAI22_X1 port map( A1 => n9007, A2 => n30385, B1 => n9775, B2 => 
                           n30379, ZN => n26556);
   U22410 : AOI221_X1 port map( B1 => n30397, B2 => n29693, C1 => n30391, C2 =>
                           n29501, A => n26530, ZN => n26521);
   U22411 : OAI22_X1 port map( A1 => n9002, A2 => n30385, B1 => n9770, B2 => 
                           n30379, ZN => n26530);
   U22412 : AOI221_X1 port map( B1 => n30397, B2 => n29694, C1 => n30391, C2 =>
                           n29502, A => n26504, ZN => n26495);
   U22413 : OAI22_X1 port map( A1 => n8997, A2 => n30385, B1 => n9765, B2 => 
                           n30379, ZN => n26504);
   U22414 : AOI221_X1 port map( B1 => n30397, B2 => n29695, C1 => n30391, C2 =>
                           n29503, A => n26478, ZN => n26469);
   U22415 : OAI22_X1 port map( A1 => n8992, A2 => n30385, B1 => n9760, B2 => 
                           n30379, ZN => n26478);
   U22416 : AOI221_X1 port map( B1 => n30398, B2 => n29696, C1 => n30392, C2 =>
                           n29504, A => n26452, ZN => n26443);
   U22417 : OAI22_X1 port map( A1 => n8987, A2 => n30386, B1 => n9755, B2 => 
                           n30380, ZN => n26452);
   U22418 : AOI221_X1 port map( B1 => n30398, B2 => n29697, C1 => n30392, C2 =>
                           n29505, A => n26426, ZN => n26417);
   U22419 : OAI22_X1 port map( A1 => n8982, A2 => n30386, B1 => n9750, B2 => 
                           n30380, ZN => n26426);
   U22420 : AOI221_X1 port map( B1 => n30398, B2 => n29698, C1 => n30392, C2 =>
                           n29506, A => n26400, ZN => n26391);
   U22421 : OAI22_X1 port map( A1 => n8977, A2 => n30386, B1 => n9745, B2 => 
                           n30380, ZN => n26400);
   U22422 : AOI221_X1 port map( B1 => n30398, B2 => n29699, C1 => n30392, C2 =>
                           n29507, A => n26368, ZN => n26349);
   U22423 : OAI22_X1 port map( A1 => n8972, A2 => n30386, B1 => n9740, B2 => 
                           n30380, ZN => n26368);
   U22424 : AOI221_X1 port map( B1 => n30261, B2 => n21927, C1 => n30255, C2 =>
                           n9606, A => n29292, ZN => n29276);
   U22425 : OAI22_X1 port map( A1 => n9286, A2 => n30249, B1 => n25667, B2 => 
                           n30243, ZN => n29292);
   U22426 : AOI221_X1 port map( B1 => n30261, B2 => n21928, C1 => n30255, C2 =>
                           n9601, A => n29263, ZN => n29256);
   U22427 : OAI22_X1 port map( A1 => n9281, A2 => n30249, B1 => n25666, B2 => 
                           n30243, ZN => n29263);
   U22428 : AOI221_X1 port map( B1 => n30261, B2 => n21929, C1 => n30255, C2 =>
                           n9596, A => n29244, ZN => n29237);
   U22429 : OAI22_X1 port map( A1 => n9276, A2 => n30249, B1 => n25665, B2 => 
                           n30243, ZN => n29244);
   U22430 : AOI221_X1 port map( B1 => n30261, B2 => n21930, C1 => n30255, C2 =>
                           n9591, A => n29225, ZN => n29218);
   U22431 : OAI22_X1 port map( A1 => n9271, A2 => n30249, B1 => n25664, B2 => 
                           n30243, ZN => n29225);
   U22432 : AOI221_X1 port map( B1 => n30261, B2 => n21931, C1 => n30255, C2 =>
                           n9586, A => n29206, ZN => n29199);
   U22433 : OAI22_X1 port map( A1 => n9266, A2 => n30249, B1 => n25663, B2 => 
                           n30243, ZN => n29206);
   U22434 : AOI221_X1 port map( B1 => n30261, B2 => n21932, C1 => n30255, C2 =>
                           n9581, A => n29187, ZN => n29180);
   U22435 : OAI22_X1 port map( A1 => n9261, A2 => n30249, B1 => n25662, B2 => 
                           n30243, ZN => n29187);
   U22436 : AOI221_X1 port map( B1 => n30261, B2 => n21933, C1 => n30255, C2 =>
                           n9576, A => n29168, ZN => n29161);
   U22437 : OAI22_X1 port map( A1 => n9256, A2 => n30249, B1 => n25661, B2 => 
                           n30243, ZN => n29168);
   U22438 : AOI221_X1 port map( B1 => n30261, B2 => n21934, C1 => n30255, C2 =>
                           n9571, A => n29149, ZN => n29142);
   U22439 : OAI22_X1 port map( A1 => n9251, A2 => n30249, B1 => n25660, B2 => 
                           n30243, ZN => n29149);
   U22440 : AOI221_X1 port map( B1 => n30261, B2 => n21935, C1 => n30255, C2 =>
                           n9566, A => n29130, ZN => n29123);
   U22441 : OAI22_X1 port map( A1 => n9246, A2 => n30249, B1 => n25659, B2 => 
                           n30243, ZN => n29130);
   U22442 : AOI221_X1 port map( B1 => n30261, B2 => n21936, C1 => n30255, C2 =>
                           n9561, A => n29111, ZN => n29104);
   U22443 : OAI22_X1 port map( A1 => n9241, A2 => n30249, B1 => n25658, B2 => 
                           n30243, ZN => n29111);
   U22444 : AOI221_X1 port map( B1 => n30261, B2 => n21937, C1 => n30255, C2 =>
                           n9556, A => n29092, ZN => n29085);
   U22445 : OAI22_X1 port map( A1 => n9236, A2 => n30249, B1 => n25657, B2 => 
                           n30243, ZN => n29092);
   U22446 : AOI221_X1 port map( B1 => n30261, B2 => n21938, C1 => n30255, C2 =>
                           n9551, A => n29073, ZN => n29066);
   U22447 : OAI22_X1 port map( A1 => n9231, A2 => n30249, B1 => n9999, B2 => 
                           n30243, ZN => n29073);
   U22448 : AOI221_X1 port map( B1 => n30262, B2 => n21939, C1 => n30256, C2 =>
                           n9546, A => n29054, ZN => n29047);
   U22449 : OAI22_X1 port map( A1 => n9226, A2 => n30250, B1 => n9994, B2 => 
                           n30244, ZN => n29054);
   U22450 : AOI221_X1 port map( B1 => n30262, B2 => n21940, C1 => n30256, C2 =>
                           n9541, A => n29035, ZN => n29028);
   U22451 : OAI22_X1 port map( A1 => n9221, A2 => n30250, B1 => n9989, B2 => 
                           n30244, ZN => n29035);
   U22452 : AOI221_X1 port map( B1 => n30262, B2 => n21941, C1 => n30256, C2 =>
                           n9536, A => n29016, ZN => n29009);
   U22453 : OAI22_X1 port map( A1 => n9216, A2 => n30250, B1 => n9984, B2 => 
                           n30244, ZN => n29016);
   U22454 : AOI221_X1 port map( B1 => n30262, B2 => n21942, C1 => n30256, C2 =>
                           n9531, A => n28997, ZN => n28990);
   U22455 : OAI22_X1 port map( A1 => n9211, A2 => n30250, B1 => n9979, B2 => 
                           n30244, ZN => n28997);
   U22456 : AOI221_X1 port map( B1 => n30262, B2 => n21943, C1 => n30256, C2 =>
                           n9526, A => n28978, ZN => n28971);
   U22457 : OAI22_X1 port map( A1 => n9206, A2 => n30250, B1 => n9974, B2 => 
                           n30244, ZN => n28978);
   U22458 : AOI221_X1 port map( B1 => n30262, B2 => n21944, C1 => n30256, C2 =>
                           n9521, A => n28959, ZN => n28952);
   U22459 : OAI22_X1 port map( A1 => n9201, A2 => n30250, B1 => n9969, B2 => 
                           n30244, ZN => n28959);
   U22460 : AOI221_X1 port map( B1 => n30262, B2 => n21945, C1 => n30256, C2 =>
                           n9516, A => n28940, ZN => n28933);
   U22461 : OAI22_X1 port map( A1 => n9196, A2 => n30250, B1 => n9964, B2 => 
                           n30244, ZN => n28940);
   U22462 : AOI221_X1 port map( B1 => n30262, B2 => n21946, C1 => n30256, C2 =>
                           n9511, A => n28921, ZN => n28914);
   U22463 : OAI22_X1 port map( A1 => n9191, A2 => n30250, B1 => n9959, B2 => 
                           n30244, ZN => n28921);
   U22464 : AOI221_X1 port map( B1 => n30262, B2 => n21947, C1 => n30256, C2 =>
                           n9506, A => n28902, ZN => n28895);
   U22465 : OAI22_X1 port map( A1 => n9186, A2 => n30250, B1 => n9954, B2 => 
                           n30244, ZN => n28902);
   U22466 : AOI221_X1 port map( B1 => n30262, B2 => n21948, C1 => n30256, C2 =>
                           n9501, A => n28883, ZN => n28876);
   U22467 : OAI22_X1 port map( A1 => n9181, A2 => n30250, B1 => n9949, B2 => 
                           n30244, ZN => n28883);
   U22468 : AOI221_X1 port map( B1 => n30262, B2 => n21949, C1 => n30256, C2 =>
                           n9496, A => n28864, ZN => n28857);
   U22469 : OAI22_X1 port map( A1 => n9176, A2 => n30250, B1 => n9944, B2 => 
                           n30244, ZN => n28864);
   U22470 : AOI221_X1 port map( B1 => n30262, B2 => n21950, C1 => n30256, C2 =>
                           n9491, A => n28845, ZN => n28838);
   U22471 : OAI22_X1 port map( A1 => n9171, A2 => n30250, B1 => n9939, B2 => 
                           n30244, ZN => n28845);
   U22472 : AOI221_X1 port map( B1 => n30263, B2 => n21951, C1 => n30257, C2 =>
                           n9486, A => n28826, ZN => n28819);
   U22473 : OAI22_X1 port map( A1 => n9166, A2 => n30251, B1 => n9934, B2 => 
                           n30245, ZN => n28826);
   U22474 : AOI221_X1 port map( B1 => n30263, B2 => n21952, C1 => n30257, C2 =>
                           n9481, A => n28807, ZN => n28800);
   U22475 : OAI22_X1 port map( A1 => n9161, A2 => n30251, B1 => n9929, B2 => 
                           n30245, ZN => n28807);
   U22476 : AOI221_X1 port map( B1 => n30263, B2 => n21953, C1 => n30257, C2 =>
                           n9476, A => n28788, ZN => n28781);
   U22477 : OAI22_X1 port map( A1 => n9156, A2 => n30251, B1 => n9924, B2 => 
                           n30245, ZN => n28788);
   U22478 : AOI221_X1 port map( B1 => n30263, B2 => n21954, C1 => n30257, C2 =>
                           n9471, A => n28769, ZN => n28762);
   U22479 : OAI22_X1 port map( A1 => n9151, A2 => n30251, B1 => n9919, B2 => 
                           n30245, ZN => n28769);
   U22480 : AOI221_X1 port map( B1 => n30263, B2 => n21955, C1 => n30257, C2 =>
                           n9466, A => n28750, ZN => n28743);
   U22481 : OAI22_X1 port map( A1 => n9146, A2 => n30251, B1 => n9914, B2 => 
                           n30245, ZN => n28750);
   U22482 : AOI221_X1 port map( B1 => n30263, B2 => n21956, C1 => n30257, C2 =>
                           n9461, A => n28731, ZN => n28724);
   U22483 : OAI22_X1 port map( A1 => n9141, A2 => n30251, B1 => n9909, B2 => 
                           n30245, ZN => n28731);
   U22484 : AOI221_X1 port map( B1 => n30263, B2 => n21957, C1 => n30257, C2 =>
                           n9456, A => n28712, ZN => n28705);
   U22485 : OAI22_X1 port map( A1 => n9136, A2 => n30251, B1 => n9904, B2 => 
                           n30245, ZN => n28712);
   U22486 : AOI221_X1 port map( B1 => n30263, B2 => n21958, C1 => n30257, C2 =>
                           n9451, A => n28693, ZN => n28686);
   U22487 : OAI22_X1 port map( A1 => n9131, A2 => n30251, B1 => n9899, B2 => 
                           n30245, ZN => n28693);
   U22488 : AOI221_X1 port map( B1 => n30263, B2 => n21959, C1 => n30257, C2 =>
                           n9446, A => n28674, ZN => n28667);
   U22489 : OAI22_X1 port map( A1 => n9126, A2 => n30251, B1 => n9894, B2 => 
                           n30245, ZN => n28674);
   U22490 : AOI221_X1 port map( B1 => n30263, B2 => n21960, C1 => n30257, C2 =>
                           n9441, A => n28655, ZN => n28648);
   U22491 : OAI22_X1 port map( A1 => n9121, A2 => n30251, B1 => n9889, B2 => 
                           n30245, ZN => n28655);
   U22492 : AOI221_X1 port map( B1 => n30263, B2 => n21961, C1 => n30257, C2 =>
                           n9436, A => n28636, ZN => n28629);
   U22493 : OAI22_X1 port map( A1 => n9116, A2 => n30251, B1 => n9884, B2 => 
                           n30245, ZN => n28636);
   U22494 : AOI221_X1 port map( B1 => n30263, B2 => n21962, C1 => n30257, C2 =>
                           n9431, A => n28617, ZN => n28610);
   U22495 : OAI22_X1 port map( A1 => n9111, A2 => n30251, B1 => n9879, B2 => 
                           n30245, ZN => n28617);
   U22496 : AOI221_X1 port map( B1 => n30264, B2 => n21963, C1 => n30258, C2 =>
                           n9426, A => n28598, ZN => n28591);
   U22497 : OAI22_X1 port map( A1 => n9106, A2 => n30252, B1 => n9874, B2 => 
                           n30246, ZN => n28598);
   U22498 : AOI221_X1 port map( B1 => n30264, B2 => n21964, C1 => n30258, C2 =>
                           n9421, A => n28579, ZN => n28572);
   U22499 : OAI22_X1 port map( A1 => n9101, A2 => n30252, B1 => n9869, B2 => 
                           n30246, ZN => n28579);
   U22500 : AOI221_X1 port map( B1 => n30264, B2 => n21965, C1 => n30258, C2 =>
                           n9416, A => n28560, ZN => n28553);
   U22501 : OAI22_X1 port map( A1 => n9096, A2 => n30252, B1 => n9864, B2 => 
                           n30246, ZN => n28560);
   U22502 : AOI221_X1 port map( B1 => n30264, B2 => n21966, C1 => n30258, C2 =>
                           n9411, A => n28541, ZN => n28534);
   U22503 : OAI22_X1 port map( A1 => n9091, A2 => n30252, B1 => n9859, B2 => 
                           n30246, ZN => n28541);
   U22504 : AOI221_X1 port map( B1 => n30264, B2 => n21967, C1 => n30258, C2 =>
                           n9406, A => n28522, ZN => n28515);
   U22505 : OAI22_X1 port map( A1 => n9086, A2 => n30252, B1 => n9854, B2 => 
                           n30246, ZN => n28522);
   U22506 : AOI221_X1 port map( B1 => n30264, B2 => n21968, C1 => n30258, C2 =>
                           n9401, A => n28503, ZN => n28496);
   U22507 : OAI22_X1 port map( A1 => n9081, A2 => n30252, B1 => n9849, B2 => 
                           n30246, ZN => n28503);
   U22508 : AOI221_X1 port map( B1 => n30264, B2 => n21969, C1 => n30258, C2 =>
                           n9396, A => n28484, ZN => n28477);
   U22509 : OAI22_X1 port map( A1 => n9076, A2 => n30252, B1 => n9844, B2 => 
                           n30246, ZN => n28484);
   U22510 : AOI221_X1 port map( B1 => n30264, B2 => n21970, C1 => n30258, C2 =>
                           n9391, A => n28465, ZN => n28458);
   U22511 : OAI22_X1 port map( A1 => n9071, A2 => n30252, B1 => n9839, B2 => 
                           n30246, ZN => n28465);
   U22512 : AOI221_X1 port map( B1 => n30264, B2 => n21971, C1 => n30258, C2 =>
                           n9386, A => n28446, ZN => n28439);
   U22513 : OAI22_X1 port map( A1 => n9066, A2 => n30252, B1 => n9834, B2 => 
                           n30246, ZN => n28446);
   U22514 : AOI221_X1 port map( B1 => n30264, B2 => n21972, C1 => n30258, C2 =>
                           n9381, A => n28427, ZN => n28420);
   U22515 : OAI22_X1 port map( A1 => n9061, A2 => n30252, B1 => n9829, B2 => 
                           n30246, ZN => n28427);
   U22516 : AOI221_X1 port map( B1 => n30264, B2 => n21973, C1 => n30258, C2 =>
                           n9376, A => n28408, ZN => n28401);
   U22517 : OAI22_X1 port map( A1 => n9056, A2 => n30252, B1 => n9824, B2 => 
                           n30246, ZN => n28408);
   U22518 : AOI221_X1 port map( B1 => n30264, B2 => n21974, C1 => n30258, C2 =>
                           n9371, A => n28389, ZN => n28382);
   U22519 : OAI22_X1 port map( A1 => n9051, A2 => n30252, B1 => n9819, B2 => 
                           n30246, ZN => n28389);
   U22520 : AOI221_X1 port map( B1 => n30265, B2 => n21975, C1 => n30259, C2 =>
                           n9366, A => n28370, ZN => n28363);
   U22521 : OAI22_X1 port map( A1 => n9046, A2 => n30253, B1 => n9814, B2 => 
                           n30247, ZN => n28370);
   U22522 : AOI221_X1 port map( B1 => n30265, B2 => n21976, C1 => n30259, C2 =>
                           n9361, A => n28351, ZN => n28344);
   U22523 : OAI22_X1 port map( A1 => n9041, A2 => n30253, B1 => n9809, B2 => 
                           n30247, ZN => n28351);
   U22524 : AOI221_X1 port map( B1 => n30265, B2 => n21977, C1 => n30259, C2 =>
                           n9356, A => n28332, ZN => n28325);
   U22525 : OAI22_X1 port map( A1 => n9036, A2 => n30253, B1 => n9804, B2 => 
                           n30247, ZN => n28332);
   U22526 : AOI221_X1 port map( B1 => n30265, B2 => n21978, C1 => n30259, C2 =>
                           n9351, A => n28313, ZN => n28306);
   U22527 : OAI22_X1 port map( A1 => n9031, A2 => n30253, B1 => n9799, B2 => 
                           n30247, ZN => n28313);
   U22528 : AOI221_X1 port map( B1 => n30265, B2 => n21979, C1 => n30259, C2 =>
                           n9346, A => n28294, ZN => n28287);
   U22529 : OAI22_X1 port map( A1 => n9026, A2 => n30253, B1 => n9794, B2 => 
                           n30247, ZN => n28294);
   U22530 : AOI221_X1 port map( B1 => n30265, B2 => n21980, C1 => n30259, C2 =>
                           n9341, A => n28275, ZN => n28268);
   U22531 : OAI22_X1 port map( A1 => n9021, A2 => n30253, B1 => n9789, B2 => 
                           n30247, ZN => n28275);
   U22532 : AOI221_X1 port map( B1 => n30265, B2 => n21981, C1 => n30259, C2 =>
                           n9336, A => n28256, ZN => n28249);
   U22533 : OAI22_X1 port map( A1 => n9016, A2 => n30253, B1 => n9784, B2 => 
                           n30247, ZN => n28256);
   U22534 : AOI221_X1 port map( B1 => n30265, B2 => n21982, C1 => n30259, C2 =>
                           n9331, A => n28237, ZN => n28230);
   U22535 : OAI22_X1 port map( A1 => n9011, A2 => n30253, B1 => n9779, B2 => 
                           n30247, ZN => n28237);
   U22536 : AOI221_X1 port map( B1 => n30265, B2 => n21983, C1 => n30259, C2 =>
                           n9326, A => n28218, ZN => n28211);
   U22537 : OAI22_X1 port map( A1 => n9006, A2 => n30253, B1 => n9774, B2 => 
                           n30247, ZN => n28218);
   U22538 : AOI221_X1 port map( B1 => n30265, B2 => n21984, C1 => n30259, C2 =>
                           n9321, A => n28199, ZN => n28192);
   U22539 : OAI22_X1 port map( A1 => n9001, A2 => n30253, B1 => n9769, B2 => 
                           n30247, ZN => n28199);
   U22540 : AOI221_X1 port map( B1 => n30265, B2 => n21985, C1 => n30259, C2 =>
                           n9316, A => n28180, ZN => n28173);
   U22541 : OAI22_X1 port map( A1 => n8996, A2 => n30253, B1 => n9764, B2 => 
                           n30247, ZN => n28180);
   U22542 : AOI221_X1 port map( B1 => n30265, B2 => n21986, C1 => n30259, C2 =>
                           n9311, A => n28161, ZN => n28154);
   U22543 : OAI22_X1 port map( A1 => n8991, A2 => n30253, B1 => n9759, B2 => 
                           n30247, ZN => n28161);
   U22544 : AOI221_X1 port map( B1 => n30266, B2 => n22012, C1 => n30260, C2 =>
                           n9306, A => n28142, ZN => n28135);
   U22545 : OAI22_X1 port map( A1 => n8986, A2 => n30254, B1 => n9754, B2 => 
                           n30248, ZN => n28142);
   U22546 : AOI221_X1 port map( B1 => n30266, B2 => n22013, C1 => n30260, C2 =>
                           n9301, A => n28123, ZN => n28116);
   U22547 : OAI22_X1 port map( A1 => n8981, A2 => n30254, B1 => n9749, B2 => 
                           n30248, ZN => n28123);
   U22548 : AOI221_X1 port map( B1 => n30266, B2 => n22014, C1 => n30260, C2 =>
                           n9296, A => n28104, ZN => n28097);
   U22549 : OAI22_X1 port map( A1 => n8976, A2 => n30254, B1 => n9744, B2 => 
                           n30248, ZN => n28104);
   U22550 : AOI221_X1 port map( B1 => n30266, B2 => n22015, C1 => n30260, C2 =>
                           n9291, A => n28066, ZN => n28045);
   U22551 : OAI22_X1 port map( A1 => n8971, A2 => n30254, B1 => n9739, B2 => 
                           n30248, ZN => n28066);
   U22552 : AOI221_X1 port map( B1 => n30466, B2 => n21987, C1 => n30460, C2 =>
                           n9607, A => n28011, ZN => n27995);
   U22553 : OAI22_X1 port map( A1 => n30459, A2 => n27990, B1 => n26315, B2 => 
                           n30447, ZN => n28011);
   U22554 : AOI221_X1 port map( B1 => n30466, B2 => n21988, C1 => n30460, C2 =>
                           n9602, A => n27975, ZN => n27968);
   U22555 : OAI22_X1 port map( A1 => n30459, A2 => n27964, B1 => n26314, B2 => 
                           n30447, ZN => n27975);
   U22556 : AOI221_X1 port map( B1 => n30466, B2 => n21989, C1 => n30460, C2 =>
                           n9597, A => n27949, ZN => n27942);
   U22557 : OAI22_X1 port map( A1 => n30459, A2 => n27938, B1 => n26313, B2 => 
                           n30447, ZN => n27949);
   U22558 : AOI221_X1 port map( B1 => n30466, B2 => n21990, C1 => n30460, C2 =>
                           n9592, A => n27923, ZN => n27916);
   U22559 : OAI22_X1 port map( A1 => n30459, A2 => n27912, B1 => n26312, B2 => 
                           n30447, ZN => n27923);
   U22560 : AOI221_X1 port map( B1 => n30466, B2 => n21991, C1 => n30460, C2 =>
                           n9587, A => n27897, ZN => n27890);
   U22561 : OAI22_X1 port map( A1 => n30459, A2 => n27886, B1 => n26311, B2 => 
                           n30447, ZN => n27897);
   U22562 : AOI221_X1 port map( B1 => n30466, B2 => n21992, C1 => n30460, C2 =>
                           n9582, A => n27871, ZN => n27864);
   U22563 : OAI22_X1 port map( A1 => n30459, A2 => n27860, B1 => n26310, B2 => 
                           n30447, ZN => n27871);
   U22564 : AOI221_X1 port map( B1 => n30466, B2 => n21993, C1 => n30460, C2 =>
                           n9577, A => n27845, ZN => n27838);
   U22565 : OAI22_X1 port map( A1 => n30459, A2 => n27834, B1 => n26309, B2 => 
                           n30447, ZN => n27845);
   U22566 : AOI221_X1 port map( B1 => n30466, B2 => n21994, C1 => n30460, C2 =>
                           n9572, A => n27819, ZN => n27812);
   U22567 : OAI22_X1 port map( A1 => n30459, A2 => n27808, B1 => n26308, B2 => 
                           n30447, ZN => n27819);
   U22568 : AOI221_X1 port map( B1 => n30466, B2 => n21995, C1 => n30460, C2 =>
                           n9567, A => n27793, ZN => n27786);
   U22569 : OAI22_X1 port map( A1 => n30459, A2 => n27782, B1 => n26307, B2 => 
                           n30447, ZN => n27793);
   U22570 : AOI221_X1 port map( B1 => n30466, B2 => n21996, C1 => n30460, C2 =>
                           n9562, A => n27767, ZN => n27760);
   U22571 : OAI22_X1 port map( A1 => n30459, A2 => n27756, B1 => n26306, B2 => 
                           n30447, ZN => n27767);
   U22572 : AOI221_X1 port map( B1 => n30466, B2 => n21997, C1 => n30460, C2 =>
                           n9557, A => n27741, ZN => n27734);
   U22573 : OAI22_X1 port map( A1 => n30459, A2 => n27730, B1 => n26305, B2 => 
                           n30447, ZN => n27741);
   U22574 : AOI221_X1 port map( B1 => n30466, B2 => n21998, C1 => n30460, C2 =>
                           n9552, A => n27715, ZN => n27708);
   U22575 : OAI22_X1 port map( A1 => n30459, A2 => n27704, B1 => n26304, B2 => 
                           n30447, ZN => n27715);
   U22576 : AOI221_X1 port map( B1 => n30467, B2 => n22076, C1 => n30461, C2 =>
                           n9547, A => n27689, ZN => n27682);
   U22577 : OAI22_X1 port map( A1 => n30458, A2 => n27678, B1 => n26303, B2 => 
                           n30448, ZN => n27689);
   U22578 : AOI221_X1 port map( B1 => n30467, B2 => n22077, C1 => n30461, C2 =>
                           n9542, A => n27663, ZN => n27656);
   U22579 : OAI22_X1 port map( A1 => n30458, A2 => n27652, B1 => n26302, B2 => 
                           n30448, ZN => n27663);
   U22580 : AOI221_X1 port map( B1 => n30467, B2 => n22078, C1 => n30461, C2 =>
                           n9537, A => n27637, ZN => n27630);
   U22581 : OAI22_X1 port map( A1 => n30458, A2 => n27626, B1 => n26301, B2 => 
                           n30448, ZN => n27637);
   U22582 : AOI221_X1 port map( B1 => n30467, B2 => n22079, C1 => n30461, C2 =>
                           n9532, A => n27611, ZN => n27604);
   U22583 : OAI22_X1 port map( A1 => n30458, A2 => n27600, B1 => n26300, B2 => 
                           n30448, ZN => n27611);
   U22584 : AOI221_X1 port map( B1 => n30467, B2 => n22080, C1 => n30461, C2 =>
                           n9527, A => n27585, ZN => n27578);
   U22585 : OAI22_X1 port map( A1 => n30458, A2 => n27574, B1 => n26299, B2 => 
                           n30448, ZN => n27585);
   U22586 : AOI221_X1 port map( B1 => n30467, B2 => n22081, C1 => n30461, C2 =>
                           n9522, A => n27559, ZN => n27552);
   U22587 : OAI22_X1 port map( A1 => n30458, A2 => n27548, B1 => n26298, B2 => 
                           n30448, ZN => n27559);
   U22588 : AOI221_X1 port map( B1 => n30467, B2 => n22082, C1 => n30461, C2 =>
                           n9517, A => n27533, ZN => n27526);
   U22589 : OAI22_X1 port map( A1 => n30458, A2 => n27522, B1 => n26297, B2 => 
                           n30448, ZN => n27533);
   U22590 : AOI221_X1 port map( B1 => n30467, B2 => n22083, C1 => n30461, C2 =>
                           n9512, A => n27507, ZN => n27500);
   U22591 : OAI22_X1 port map( A1 => n30458, A2 => n27496, B1 => n26296, B2 => 
                           n30448, ZN => n27507);
   U22592 : AOI221_X1 port map( B1 => n30467, B2 => n22084, C1 => n30461, C2 =>
                           n9507, A => n27481, ZN => n27474);
   U22593 : OAI22_X1 port map( A1 => n30458, A2 => n27470, B1 => n26295, B2 => 
                           n30448, ZN => n27481);
   U22594 : AOI221_X1 port map( B1 => n30467, B2 => n22085, C1 => n30461, C2 =>
                           n9502, A => n27455, ZN => n27448);
   U22595 : OAI22_X1 port map( A1 => n30458, A2 => n27444, B1 => n26294, B2 => 
                           n30448, ZN => n27455);
   U22596 : AOI221_X1 port map( B1 => n30467, B2 => n22086, C1 => n30461, C2 =>
                           n9497, A => n27429, ZN => n27422);
   U22597 : OAI22_X1 port map( A1 => n30458, A2 => n27418, B1 => n26293, B2 => 
                           n30448, ZN => n27429);
   U22598 : AOI221_X1 port map( B1 => n30467, B2 => n22087, C1 => n30461, C2 =>
                           n9492, A => n27403, ZN => n27396);
   U22599 : OAI22_X1 port map( A1 => n30458, A2 => n27392, B1 => n26292, B2 => 
                           n30448, ZN => n27403);
   U22600 : AOI221_X1 port map( B1 => n30468, B2 => n22088, C1 => n30462, C2 =>
                           n9487, A => n27377, ZN => n27370);
   U22601 : OAI22_X1 port map( A1 => n30458, A2 => n27366, B1 => n26291, B2 => 
                           n30449, ZN => n27377);
   U22602 : AOI221_X1 port map( B1 => n30470, B2 => n21999, C1 => n30464, C2 =>
                           n9352, A => n26675, ZN => n26668);
   U22603 : OAI22_X1 port map( A1 => n30455, A2 => n26664, B1 => n26264, B2 => 
                           n30451, ZN => n26675);
   U22604 : AOI221_X1 port map( B1 => n30470, B2 => n22000, C1 => n30464, C2 =>
                           n9347, A => n26649, ZN => n26642);
   U22605 : OAI22_X1 port map( A1 => n30455, A2 => n26638, B1 => n26263, B2 => 
                           n30451, ZN => n26649);
   U22606 : AOI221_X1 port map( B1 => n30470, B2 => n22001, C1 => n30464, C2 =>
                           n9342, A => n26623, ZN => n26616);
   U22607 : OAI22_X1 port map( A1 => n30455, A2 => n26612, B1 => n26262, B2 => 
                           n30451, ZN => n26623);
   U22608 : AOI221_X1 port map( B1 => n30470, B2 => n22002, C1 => n30464, C2 =>
                           n9337, A => n26597, ZN => n26590);
   U22609 : OAI22_X1 port map( A1 => n30455, A2 => n26586, B1 => n26261, B2 => 
                           n30451, ZN => n26597);
   U22610 : AOI221_X1 port map( B1 => n30470, B2 => n22003, C1 => n30464, C2 =>
                           n9332, A => n26571, ZN => n26564);
   U22611 : OAI22_X1 port map( A1 => n30455, A2 => n26560, B1 => n26260, B2 => 
                           n30451, ZN => n26571);
   U22612 : AOI221_X1 port map( B1 => n30470, B2 => n22004, C1 => n30464, C2 =>
                           n9327, A => n26545, ZN => n26538);
   U22613 : OAI22_X1 port map( A1 => n30455, A2 => n26534, B1 => n26259, B2 => 
                           n30451, ZN => n26545);
   U22614 : AOI221_X1 port map( B1 => n30470, B2 => n22005, C1 => n30464, C2 =>
                           n9322, A => n26519, ZN => n26512);
   U22615 : OAI22_X1 port map( A1 => n30455, A2 => n26508, B1 => n26258, B2 => 
                           n30451, ZN => n26519);
   U22616 : AOI221_X1 port map( B1 => n30470, B2 => n22006, C1 => n30464, C2 =>
                           n9317, A => n26493, ZN => n26486);
   U22617 : OAI22_X1 port map( A1 => n30455, A2 => n26482, B1 => n26257, B2 => 
                           n30451, ZN => n26493);
   U22618 : AOI221_X1 port map( B1 => n30470, B2 => n22007, C1 => n30464, C2 =>
                           n9312, A => n26467, ZN => n26460);
   U22619 : OAI22_X1 port map( A1 => n30455, A2 => n26456, B1 => n26256, B2 => 
                           n30451, ZN => n26467);
   U22620 : AOI221_X1 port map( B1 => n30471, B2 => n22008, C1 => n30465, C2 =>
                           n9307, A => n26441, ZN => n26434);
   U22621 : OAI22_X1 port map( A1 => n30455, A2 => n26430, B1 => n26255, B2 => 
                           n30452, ZN => n26441);
   U22622 : AOI221_X1 port map( B1 => n30471, B2 => n22009, C1 => n30465, C2 =>
                           n9302, A => n26415, ZN => n26408);
   U22623 : OAI22_X1 port map( A1 => n30455, A2 => n26404, B1 => n26254, B2 => 
                           n30452, ZN => n26415);
   U22624 : AOI221_X1 port map( B1 => n30471, B2 => n22010, C1 => n30465, C2 =>
                           n9297, A => n26389, ZN => n26382);
   U22625 : OAI22_X1 port map( A1 => n30455, A2 => n26378, B1 => n26253, B2 => 
                           n30452, ZN => n26389);
   U22626 : AOI221_X1 port map( B1 => n30471, B2 => n22011, C1 => n30465, C2 =>
                           n9292, A => n26345, ZN => n26324);
   U22627 : OAI22_X1 port map( A1 => n26317, A2 => n30455, B1 => n26251, B2 => 
                           n30452, ZN => n26345);
   U22628 : AOI221_X1 port map( B1 => n30165, B2 => n29700, C1 => n30159, C2 =>
                           n29508, A => n29307, ZN => n29294);
   U22629 : OAI22_X1 port map( A1 => n9288, A2 => n30153, B1 => n25954, B2 => 
                           n30147, ZN => n29307);
   U22630 : AOI221_X1 port map( B1 => n30165, B2 => n29701, C1 => n30159, C2 =>
                           n29509, A => n29271, ZN => n29264);
   U22631 : OAI22_X1 port map( A1 => n9283, A2 => n30153, B1 => n25953, B2 => 
                           n30147, ZN => n29271);
   U22632 : AOI221_X1 port map( B1 => n30165, B2 => n29702, C1 => n30159, C2 =>
                           n29510, A => n29252, ZN => n29245);
   U22633 : OAI22_X1 port map( A1 => n9278, A2 => n30153, B1 => n25952, B2 => 
                           n30147, ZN => n29252);
   U22634 : AOI221_X1 port map( B1 => n30165, B2 => n29703, C1 => n30159, C2 =>
                           n29511, A => n29233, ZN => n29226);
   U22635 : OAI22_X1 port map( A1 => n9273, A2 => n30153, B1 => n25951, B2 => 
                           n30147, ZN => n29233);
   U22636 : AOI221_X1 port map( B1 => n30165, B2 => n29704, C1 => n30159, C2 =>
                           n29512, A => n29214, ZN => n29207);
   U22637 : OAI22_X1 port map( A1 => n9268, A2 => n30153, B1 => n25950, B2 => 
                           n30147, ZN => n29214);
   U22638 : AOI221_X1 port map( B1 => n30165, B2 => n29705, C1 => n30159, C2 =>
                           n29513, A => n29195, ZN => n29188);
   U22639 : OAI22_X1 port map( A1 => n9263, A2 => n30153, B1 => n25949, B2 => 
                           n30147, ZN => n29195);
   U22640 : AOI221_X1 port map( B1 => n30165, B2 => n29706, C1 => n30159, C2 =>
                           n29514, A => n29176, ZN => n29169);
   U22641 : OAI22_X1 port map( A1 => n9258, A2 => n30153, B1 => n25948, B2 => 
                           n30147, ZN => n29176);
   U22642 : AOI221_X1 port map( B1 => n30165, B2 => n29707, C1 => n30159, C2 =>
                           n29515, A => n29157, ZN => n29150);
   U22643 : OAI22_X1 port map( A1 => n9253, A2 => n30153, B1 => n25947, B2 => 
                           n30147, ZN => n29157);
   U22644 : AOI221_X1 port map( B1 => n30165, B2 => n29708, C1 => n30159, C2 =>
                           n29516, A => n29138, ZN => n29131);
   U22645 : OAI22_X1 port map( A1 => n9248, A2 => n30153, B1 => n25946, B2 => 
                           n30147, ZN => n29138);
   U22646 : AOI221_X1 port map( B1 => n30165, B2 => n29709, C1 => n30159, C2 =>
                           n29517, A => n29119, ZN => n29112);
   U22647 : OAI22_X1 port map( A1 => n9243, A2 => n30153, B1 => n25945, B2 => 
                           n30147, ZN => n29119);
   U22648 : AOI221_X1 port map( B1 => n30165, B2 => n29710, C1 => n30159, C2 =>
                           n29518, A => n29100, ZN => n29093);
   U22649 : OAI22_X1 port map( A1 => n9238, A2 => n30153, B1 => n25944, B2 => 
                           n30147, ZN => n29100);
   U22650 : AOI221_X1 port map( B1 => n30165, B2 => n29711, C1 => n30159, C2 =>
                           n29519, A => n29081, ZN => n29074);
   U22651 : OAI22_X1 port map( A1 => n9233, A2 => n30153, B1 => n25943, B2 => 
                           n30147, ZN => n29081);
   U22652 : AOI221_X1 port map( B1 => n30166, B2 => n29712, C1 => n30160, C2 =>
                           n29520, A => n29062, ZN => n29055);
   U22653 : OAI22_X1 port map( A1 => n9228, A2 => n30154, B1 => n9996, B2 => 
                           n30148, ZN => n29062);
   U22654 : AOI221_X1 port map( B1 => n30166, B2 => n29713, C1 => n30160, C2 =>
                           n29521, A => n29043, ZN => n29036);
   U22655 : OAI22_X1 port map( A1 => n9223, A2 => n30154, B1 => n9991, B2 => 
                           n30148, ZN => n29043);
   U22656 : AOI221_X1 port map( B1 => n30166, B2 => n29714, C1 => n30160, C2 =>
                           n29522, A => n29024, ZN => n29017);
   U22657 : OAI22_X1 port map( A1 => n9218, A2 => n30154, B1 => n9986, B2 => 
                           n30148, ZN => n29024);
   U22658 : AOI221_X1 port map( B1 => n30166, B2 => n29715, C1 => n30160, C2 =>
                           n29523, A => n29005, ZN => n28998);
   U22659 : OAI22_X1 port map( A1 => n9213, A2 => n30154, B1 => n9981, B2 => 
                           n30148, ZN => n29005);
   U22660 : AOI221_X1 port map( B1 => n30166, B2 => n29716, C1 => n30160, C2 =>
                           n29524, A => n28986, ZN => n28979);
   U22661 : OAI22_X1 port map( A1 => n9208, A2 => n30154, B1 => n9976, B2 => 
                           n30148, ZN => n28986);
   U22662 : AOI221_X1 port map( B1 => n30166, B2 => n29717, C1 => n30160, C2 =>
                           n29525, A => n28967, ZN => n28960);
   U22663 : OAI22_X1 port map( A1 => n9203, A2 => n30154, B1 => n9971, B2 => 
                           n30148, ZN => n28967);
   U22664 : AOI221_X1 port map( B1 => n30166, B2 => n29718, C1 => n30160, C2 =>
                           n29526, A => n28948, ZN => n28941);
   U22665 : OAI22_X1 port map( A1 => n9198, A2 => n30154, B1 => n9966, B2 => 
                           n30148, ZN => n28948);
   U22666 : AOI221_X1 port map( B1 => n30166, B2 => n29719, C1 => n30160, C2 =>
                           n29527, A => n28929, ZN => n28922);
   U22667 : OAI22_X1 port map( A1 => n9193, A2 => n30154, B1 => n9961, B2 => 
                           n30148, ZN => n28929);
   U22668 : AOI221_X1 port map( B1 => n30166, B2 => n29720, C1 => n30160, C2 =>
                           n29528, A => n28910, ZN => n28903);
   U22669 : OAI22_X1 port map( A1 => n9188, A2 => n30154, B1 => n9956, B2 => 
                           n30148, ZN => n28910);
   U22670 : AOI221_X1 port map( B1 => n30166, B2 => n29721, C1 => n30160, C2 =>
                           n29529, A => n28891, ZN => n28884);
   U22671 : OAI22_X1 port map( A1 => n9183, A2 => n30154, B1 => n9951, B2 => 
                           n30148, ZN => n28891);
   U22672 : AOI221_X1 port map( B1 => n30166, B2 => n29722, C1 => n30160, C2 =>
                           n29530, A => n28872, ZN => n28865);
   U22673 : OAI22_X1 port map( A1 => n9178, A2 => n30154, B1 => n9946, B2 => 
                           n30148, ZN => n28872);
   U22674 : AOI221_X1 port map( B1 => n30166, B2 => n29723, C1 => n30160, C2 =>
                           n29531, A => n28853, ZN => n28846);
   U22675 : OAI22_X1 port map( A1 => n9173, A2 => n30154, B1 => n9941, B2 => 
                           n30148, ZN => n28853);
   U22676 : AOI221_X1 port map( B1 => n30167, B2 => n29724, C1 => n30161, C2 =>
                           n29532, A => n28834, ZN => n28827);
   U22677 : OAI22_X1 port map( A1 => n9168, A2 => n30155, B1 => n9936, B2 => 
                           n30149, ZN => n28834);
   U22678 : AOI221_X1 port map( B1 => n30167, B2 => n29725, C1 => n30161, C2 =>
                           n29533, A => n28815, ZN => n28808);
   U22679 : OAI22_X1 port map( A1 => n9163, A2 => n30155, B1 => n9931, B2 => 
                           n30149, ZN => n28815);
   U22680 : AOI221_X1 port map( B1 => n30167, B2 => n29726, C1 => n30161, C2 =>
                           n29534, A => n28796, ZN => n28789);
   U22681 : OAI22_X1 port map( A1 => n9158, A2 => n30155, B1 => n9926, B2 => 
                           n30149, ZN => n28796);
   U22682 : AOI221_X1 port map( B1 => n30167, B2 => n29727, C1 => n30161, C2 =>
                           n29535, A => n28777, ZN => n28770);
   U22683 : OAI22_X1 port map( A1 => n9153, A2 => n30155, B1 => n9921, B2 => 
                           n30149, ZN => n28777);
   U22684 : AOI221_X1 port map( B1 => n30167, B2 => n29728, C1 => n30161, C2 =>
                           n29536, A => n28758, ZN => n28751);
   U22685 : OAI22_X1 port map( A1 => n9148, A2 => n30155, B1 => n9916, B2 => 
                           n30149, ZN => n28758);
   U22686 : AOI221_X1 port map( B1 => n30167, B2 => n29729, C1 => n30161, C2 =>
                           n29537, A => n28739, ZN => n28732);
   U22687 : OAI22_X1 port map( A1 => n9143, A2 => n30155, B1 => n9911, B2 => 
                           n30149, ZN => n28739);
   U22688 : AOI221_X1 port map( B1 => n30167, B2 => n29730, C1 => n30161, C2 =>
                           n29538, A => n28720, ZN => n28713);
   U22689 : OAI22_X1 port map( A1 => n9138, A2 => n30155, B1 => n9906, B2 => 
                           n30149, ZN => n28720);
   U22690 : AOI221_X1 port map( B1 => n30167, B2 => n29731, C1 => n30161, C2 =>
                           n29539, A => n28701, ZN => n28694);
   U22691 : OAI22_X1 port map( A1 => n9133, A2 => n30155, B1 => n9901, B2 => 
                           n30149, ZN => n28701);
   U22692 : AOI221_X1 port map( B1 => n30167, B2 => n29732, C1 => n30161, C2 =>
                           n29540, A => n28682, ZN => n28675);
   U22693 : OAI22_X1 port map( A1 => n9128, A2 => n30155, B1 => n9896, B2 => 
                           n30149, ZN => n28682);
   U22694 : AOI221_X1 port map( B1 => n30167, B2 => n29733, C1 => n30161, C2 =>
                           n29541, A => n28663, ZN => n28656);
   U22695 : OAI22_X1 port map( A1 => n9123, A2 => n30155, B1 => n9891, B2 => 
                           n30149, ZN => n28663);
   U22696 : AOI221_X1 port map( B1 => n30167, B2 => n29734, C1 => n30161, C2 =>
                           n29542, A => n28644, ZN => n28637);
   U22697 : OAI22_X1 port map( A1 => n9118, A2 => n30155, B1 => n9886, B2 => 
                           n30149, ZN => n28644);
   U22698 : AOI221_X1 port map( B1 => n30167, B2 => n29735, C1 => n30161, C2 =>
                           n29543, A => n28625, ZN => n28618);
   U22699 : OAI22_X1 port map( A1 => n9113, A2 => n30155, B1 => n9881, B2 => 
                           n30149, ZN => n28625);
   U22700 : AOI221_X1 port map( B1 => n30168, B2 => n29736, C1 => n30162, C2 =>
                           n29544, A => n28606, ZN => n28599);
   U22701 : OAI22_X1 port map( A1 => n9108, A2 => n30156, B1 => n9876, B2 => 
                           n30150, ZN => n28606);
   U22702 : AOI221_X1 port map( B1 => n30168, B2 => n29737, C1 => n30162, C2 =>
                           n29545, A => n28587, ZN => n28580);
   U22703 : OAI22_X1 port map( A1 => n9103, A2 => n30156, B1 => n9871, B2 => 
                           n30150, ZN => n28587);
   U22704 : AOI221_X1 port map( B1 => n30168, B2 => n29738, C1 => n30162, C2 =>
                           n29546, A => n28568, ZN => n28561);
   U22705 : OAI22_X1 port map( A1 => n9098, A2 => n30156, B1 => n9866, B2 => 
                           n30150, ZN => n28568);
   U22706 : AOI221_X1 port map( B1 => n30168, B2 => n29739, C1 => n30162, C2 =>
                           n29547, A => n28549, ZN => n28542);
   U22707 : OAI22_X1 port map( A1 => n9093, A2 => n30156, B1 => n9861, B2 => 
                           n30150, ZN => n28549);
   U22708 : AOI221_X1 port map( B1 => n30168, B2 => n29740, C1 => n30162, C2 =>
                           n29548, A => n28530, ZN => n28523);
   U22709 : OAI22_X1 port map( A1 => n9088, A2 => n30156, B1 => n9856, B2 => 
                           n30150, ZN => n28530);
   U22710 : AOI221_X1 port map( B1 => n30168, B2 => n29741, C1 => n30162, C2 =>
                           n29549, A => n28511, ZN => n28504);
   U22711 : OAI22_X1 port map( A1 => n9083, A2 => n30156, B1 => n9851, B2 => 
                           n30150, ZN => n28511);
   U22712 : AOI221_X1 port map( B1 => n30168, B2 => n29742, C1 => n30162, C2 =>
                           n29550, A => n28492, ZN => n28485);
   U22713 : OAI22_X1 port map( A1 => n9078, A2 => n30156, B1 => n9846, B2 => 
                           n30150, ZN => n28492);
   U22714 : AOI221_X1 port map( B1 => n30168, B2 => n29743, C1 => n30162, C2 =>
                           n29551, A => n28473, ZN => n28466);
   U22715 : OAI22_X1 port map( A1 => n9073, A2 => n30156, B1 => n9841, B2 => 
                           n30150, ZN => n28473);
   U22716 : AOI221_X1 port map( B1 => n30168, B2 => n29744, C1 => n30162, C2 =>
                           n29552, A => n28454, ZN => n28447);
   U22717 : OAI22_X1 port map( A1 => n9068, A2 => n30156, B1 => n9836, B2 => 
                           n30150, ZN => n28454);
   U22718 : AOI221_X1 port map( B1 => n30168, B2 => n29745, C1 => n30162, C2 =>
                           n29553, A => n28435, ZN => n28428);
   U22719 : OAI22_X1 port map( A1 => n9063, A2 => n30156, B1 => n9831, B2 => 
                           n30150, ZN => n28435);
   U22720 : AOI221_X1 port map( B1 => n30168, B2 => n29746, C1 => n30162, C2 =>
                           n29554, A => n28416, ZN => n28409);
   U22721 : OAI22_X1 port map( A1 => n9058, A2 => n30156, B1 => n9826, B2 => 
                           n30150, ZN => n28416);
   U22722 : AOI221_X1 port map( B1 => n30168, B2 => n29747, C1 => n30162, C2 =>
                           n29555, A => n28397, ZN => n28390);
   U22723 : OAI22_X1 port map( A1 => n9053, A2 => n30156, B1 => n9821, B2 => 
                           n30150, ZN => n28397);
   U22724 : AOI221_X1 port map( B1 => n30169, B2 => n29748, C1 => n30163, C2 =>
                           n29556, A => n28378, ZN => n28371);
   U22725 : OAI22_X1 port map( A1 => n9048, A2 => n30157, B1 => n9816, B2 => 
                           n30151, ZN => n28378);
   U22726 : AOI221_X1 port map( B1 => n30169, B2 => n29749, C1 => n30163, C2 =>
                           n29557, A => n28359, ZN => n28352);
   U22727 : OAI22_X1 port map( A1 => n9043, A2 => n30157, B1 => n9811, B2 => 
                           n30151, ZN => n28359);
   U22728 : AOI221_X1 port map( B1 => n30169, B2 => n29750, C1 => n30163, C2 =>
                           n29558, A => n28340, ZN => n28333);
   U22729 : OAI22_X1 port map( A1 => n9038, A2 => n30157, B1 => n9806, B2 => 
                           n30151, ZN => n28340);
   U22730 : AOI221_X1 port map( B1 => n30169, B2 => n29751, C1 => n30163, C2 =>
                           n29559, A => n28321, ZN => n28314);
   U22731 : OAI22_X1 port map( A1 => n9033, A2 => n30157, B1 => n9801, B2 => 
                           n30151, ZN => n28321);
   U22732 : AOI221_X1 port map( B1 => n30169, B2 => n29752, C1 => n30163, C2 =>
                           n29560, A => n28302, ZN => n28295);
   U22733 : OAI22_X1 port map( A1 => n9028, A2 => n30157, B1 => n9796, B2 => 
                           n30151, ZN => n28302);
   U22734 : AOI221_X1 port map( B1 => n30169, B2 => n29753, C1 => n30163, C2 =>
                           n29561, A => n28283, ZN => n28276);
   U22735 : OAI22_X1 port map( A1 => n9023, A2 => n30157, B1 => n9791, B2 => 
                           n30151, ZN => n28283);
   U22736 : AOI221_X1 port map( B1 => n30169, B2 => n29754, C1 => n30163, C2 =>
                           n29562, A => n28264, ZN => n28257);
   U22737 : OAI22_X1 port map( A1 => n9018, A2 => n30157, B1 => n9786, B2 => 
                           n30151, ZN => n28264);
   U22738 : AOI221_X1 port map( B1 => n30169, B2 => n29755, C1 => n30163, C2 =>
                           n29563, A => n28245, ZN => n28238);
   U22739 : OAI22_X1 port map( A1 => n9013, A2 => n30157, B1 => n9781, B2 => 
                           n30151, ZN => n28245);
   U22740 : AOI221_X1 port map( B1 => n30169, B2 => n29756, C1 => n30163, C2 =>
                           n29564, A => n28226, ZN => n28219);
   U22741 : OAI22_X1 port map( A1 => n9008, A2 => n30157, B1 => n9776, B2 => 
                           n30151, ZN => n28226);
   U22742 : AOI221_X1 port map( B1 => n30169, B2 => n29757, C1 => n30163, C2 =>
                           n29565, A => n28207, ZN => n28200);
   U22743 : OAI22_X1 port map( A1 => n9003, A2 => n30157, B1 => n9771, B2 => 
                           n30151, ZN => n28207);
   U22744 : AOI221_X1 port map( B1 => n30169, B2 => n29758, C1 => n30163, C2 =>
                           n29566, A => n28188, ZN => n28181);
   U22745 : OAI22_X1 port map( A1 => n8998, A2 => n30157, B1 => n9766, B2 => 
                           n30151, ZN => n28188);
   U22746 : AOI221_X1 port map( B1 => n30169, B2 => n29759, C1 => n30163, C2 =>
                           n29567, A => n28169, ZN => n28162);
   U22747 : OAI22_X1 port map( A1 => n8993, A2 => n30157, B1 => n9761, B2 => 
                           n30151, ZN => n28169);
   U22748 : AOI221_X1 port map( B1 => n30170, B2 => n29760, C1 => n30164, C2 =>
                           n29568, A => n28150, ZN => n28143);
   U22749 : OAI22_X1 port map( A1 => n8988, A2 => n30158, B1 => n9756, B2 => 
                           n30152, ZN => n28150);
   U22750 : AOI221_X1 port map( B1 => n30170, B2 => n29761, C1 => n30164, C2 =>
                           n29569, A => n28131, ZN => n28124);
   U22751 : OAI22_X1 port map( A1 => n8983, A2 => n30158, B1 => n9751, B2 => 
                           n30152, ZN => n28131);
   U22752 : AOI221_X1 port map( B1 => n30170, B2 => n29762, C1 => n30164, C2 =>
                           n29570, A => n28112, ZN => n28105);
   U22753 : OAI22_X1 port map( A1 => n8978, A2 => n30158, B1 => n9746, B2 => 
                           n30152, ZN => n28112);
   U22754 : AOI221_X1 port map( B1 => n30170, B2 => n29763, C1 => n30164, C2 =>
                           n29571, A => n28090, ZN => n28069);
   U22755 : OAI22_X1 port map( A1 => n8973, A2 => n30158, B1 => n9741, B2 => 
                           n30152, ZN => n28090);
   U22756 : AOI221_X1 port map( B1 => n30369, B2 => n29700, C1 => n30363, C2 =>
                           n29508, A => n28032, ZN => n28014);
   U22757 : OAI22_X1 port map( A1 => n9288, A2 => n30357, B1 => n25954, B2 => 
                           n30351, ZN => n28032);
   U22758 : AOI221_X1 port map( B1 => n30369, B2 => n29701, C1 => n30363, C2 =>
                           n29509, A => n27989, ZN => n27976);
   U22759 : OAI22_X1 port map( A1 => n9283, A2 => n30357, B1 => n25953, B2 => 
                           n30351, ZN => n27989);
   U22760 : AOI221_X1 port map( B1 => n30369, B2 => n29702, C1 => n30363, C2 =>
                           n29510, A => n27963, ZN => n27950);
   U22761 : OAI22_X1 port map( A1 => n9278, A2 => n30357, B1 => n25952, B2 => 
                           n30351, ZN => n27963);
   U22762 : AOI221_X1 port map( B1 => n30369, B2 => n29703, C1 => n30363, C2 =>
                           n29511, A => n27937, ZN => n27924);
   U22763 : OAI22_X1 port map( A1 => n9273, A2 => n30357, B1 => n25951, B2 => 
                           n30351, ZN => n27937);
   U22764 : AOI221_X1 port map( B1 => n30369, B2 => n29704, C1 => n30363, C2 =>
                           n29512, A => n27911, ZN => n27898);
   U22765 : OAI22_X1 port map( A1 => n9268, A2 => n30357, B1 => n25950, B2 => 
                           n30351, ZN => n27911);
   U22766 : AOI221_X1 port map( B1 => n30369, B2 => n29705, C1 => n30363, C2 =>
                           n29513, A => n27885, ZN => n27872);
   U22767 : OAI22_X1 port map( A1 => n9263, A2 => n30357, B1 => n25949, B2 => 
                           n30351, ZN => n27885);
   U22768 : AOI221_X1 port map( B1 => n30369, B2 => n29706, C1 => n30363, C2 =>
                           n29514, A => n27859, ZN => n27846);
   U22769 : OAI22_X1 port map( A1 => n9258, A2 => n30357, B1 => n25948, B2 => 
                           n30351, ZN => n27859);
   U22770 : AOI221_X1 port map( B1 => n30369, B2 => n29707, C1 => n30363, C2 =>
                           n29515, A => n27833, ZN => n27820);
   U22771 : OAI22_X1 port map( A1 => n9253, A2 => n30357, B1 => n25947, B2 => 
                           n30351, ZN => n27833);
   U22772 : AOI221_X1 port map( B1 => n30369, B2 => n29708, C1 => n30363, C2 =>
                           n29516, A => n27807, ZN => n27794);
   U22773 : OAI22_X1 port map( A1 => n9248, A2 => n30357, B1 => n25946, B2 => 
                           n30351, ZN => n27807);
   U22774 : AOI221_X1 port map( B1 => n30369, B2 => n29709, C1 => n30363, C2 =>
                           n29517, A => n27781, ZN => n27768);
   U22775 : OAI22_X1 port map( A1 => n9243, A2 => n30357, B1 => n25945, B2 => 
                           n30351, ZN => n27781);
   U22776 : AOI221_X1 port map( B1 => n30369, B2 => n29710, C1 => n30363, C2 =>
                           n29518, A => n27755, ZN => n27742);
   U22777 : OAI22_X1 port map( A1 => n9238, A2 => n30357, B1 => n25944, B2 => 
                           n30351, ZN => n27755);
   U22778 : AOI221_X1 port map( B1 => n30369, B2 => n29711, C1 => n30363, C2 =>
                           n29519, A => n27729, ZN => n27716);
   U22779 : OAI22_X1 port map( A1 => n9233, A2 => n30357, B1 => n25943, B2 => 
                           n30351, ZN => n27729);
   U22780 : AOI221_X1 port map( B1 => n30370, B2 => n29712, C1 => n30364, C2 =>
                           n29520, A => n27703, ZN => n27690);
   U22781 : OAI22_X1 port map( A1 => n9228, A2 => n30358, B1 => n9996, B2 => 
                           n30352, ZN => n27703);
   U22782 : AOI221_X1 port map( B1 => n30370, B2 => n29713, C1 => n30364, C2 =>
                           n29521, A => n27677, ZN => n27664);
   U22783 : OAI22_X1 port map( A1 => n9223, A2 => n30358, B1 => n9991, B2 => 
                           n30352, ZN => n27677);
   U22784 : AOI221_X1 port map( B1 => n30370, B2 => n29714, C1 => n30364, C2 =>
                           n29522, A => n27651, ZN => n27638);
   U22785 : OAI22_X1 port map( A1 => n9218, A2 => n30358, B1 => n9986, B2 => 
                           n30352, ZN => n27651);
   U22786 : AOI221_X1 port map( B1 => n30370, B2 => n29715, C1 => n30364, C2 =>
                           n29523, A => n27625, ZN => n27612);
   U22787 : OAI22_X1 port map( A1 => n9213, A2 => n30358, B1 => n9981, B2 => 
                           n30352, ZN => n27625);
   U22788 : AOI221_X1 port map( B1 => n30370, B2 => n29716, C1 => n30364, C2 =>
                           n29524, A => n27599, ZN => n27586);
   U22789 : OAI22_X1 port map( A1 => n9208, A2 => n30358, B1 => n9976, B2 => 
                           n30352, ZN => n27599);
   U22790 : AOI221_X1 port map( B1 => n30370, B2 => n29717, C1 => n30364, C2 =>
                           n29525, A => n27573, ZN => n27560);
   U22791 : OAI22_X1 port map( A1 => n9203, A2 => n30358, B1 => n9971, B2 => 
                           n30352, ZN => n27573);
   U22792 : AOI221_X1 port map( B1 => n30370, B2 => n29718, C1 => n30364, C2 =>
                           n29526, A => n27547, ZN => n27534);
   U22793 : OAI22_X1 port map( A1 => n9198, A2 => n30358, B1 => n9966, B2 => 
                           n30352, ZN => n27547);
   U22794 : AOI221_X1 port map( B1 => n30370, B2 => n29719, C1 => n30364, C2 =>
                           n29527, A => n27521, ZN => n27508);
   U22795 : OAI22_X1 port map( A1 => n9193, A2 => n30358, B1 => n9961, B2 => 
                           n30352, ZN => n27521);
   U22796 : AOI221_X1 port map( B1 => n30370, B2 => n29720, C1 => n30364, C2 =>
                           n29528, A => n27495, ZN => n27482);
   U22797 : OAI22_X1 port map( A1 => n9188, A2 => n30358, B1 => n9956, B2 => 
                           n30352, ZN => n27495);
   U22798 : AOI221_X1 port map( B1 => n30370, B2 => n29721, C1 => n30364, C2 =>
                           n29529, A => n27469, ZN => n27456);
   U22799 : OAI22_X1 port map( A1 => n9183, A2 => n30358, B1 => n9951, B2 => 
                           n30352, ZN => n27469);
   U22800 : AOI221_X1 port map( B1 => n30370, B2 => n29722, C1 => n30364, C2 =>
                           n29530, A => n27443, ZN => n27430);
   U22801 : OAI22_X1 port map( A1 => n9178, A2 => n30358, B1 => n9946, B2 => 
                           n30352, ZN => n27443);
   U22802 : AOI221_X1 port map( B1 => n30370, B2 => n29723, C1 => n30364, C2 =>
                           n29531, A => n27417, ZN => n27404);
   U22803 : OAI22_X1 port map( A1 => n9173, A2 => n30358, B1 => n9941, B2 => 
                           n30352, ZN => n27417);
   U22804 : AOI221_X1 port map( B1 => n30371, B2 => n29724, C1 => n30365, C2 =>
                           n29532, A => n27391, ZN => n27378);
   U22805 : OAI22_X1 port map( A1 => n9168, A2 => n30359, B1 => n9936, B2 => 
                           n30353, ZN => n27391);
   U22806 : AOI221_X1 port map( B1 => n30371, B2 => n29725, C1 => n30365, C2 =>
                           n29533, A => n27365, ZN => n27352);
   U22807 : OAI22_X1 port map( A1 => n9163, A2 => n30359, B1 => n9931, B2 => 
                           n30353, ZN => n27365);
   U22808 : AOI221_X1 port map( B1 => n30371, B2 => n29726, C1 => n30365, C2 =>
                           n29534, A => n27339, ZN => n27326);
   U22809 : OAI22_X1 port map( A1 => n9158, A2 => n30359, B1 => n9926, B2 => 
                           n30353, ZN => n27339);
   U22810 : AOI221_X1 port map( B1 => n30371, B2 => n29727, C1 => n30365, C2 =>
                           n29535, A => n27313, ZN => n27300);
   U22811 : OAI22_X1 port map( A1 => n9153, A2 => n30359, B1 => n9921, B2 => 
                           n30353, ZN => n27313);
   U22812 : AOI221_X1 port map( B1 => n30371, B2 => n29728, C1 => n30365, C2 =>
                           n29536, A => n27287, ZN => n27274);
   U22813 : OAI22_X1 port map( A1 => n9148, A2 => n30359, B1 => n9916, B2 => 
                           n30353, ZN => n27287);
   U22814 : AOI221_X1 port map( B1 => n30371, B2 => n29729, C1 => n30365, C2 =>
                           n29537, A => n27261, ZN => n27248);
   U22815 : OAI22_X1 port map( A1 => n9143, A2 => n30359, B1 => n9911, B2 => 
                           n30353, ZN => n27261);
   U22816 : AOI221_X1 port map( B1 => n30371, B2 => n29730, C1 => n30365, C2 =>
                           n29538, A => n27235, ZN => n27222);
   U22817 : OAI22_X1 port map( A1 => n9138, A2 => n30359, B1 => n9906, B2 => 
                           n30353, ZN => n27235);
   U22818 : AOI221_X1 port map( B1 => n30371, B2 => n29731, C1 => n30365, C2 =>
                           n29539, A => n27209, ZN => n27196);
   U22819 : OAI22_X1 port map( A1 => n9133, A2 => n30359, B1 => n9901, B2 => 
                           n30353, ZN => n27209);
   U22820 : AOI221_X1 port map( B1 => n30371, B2 => n29732, C1 => n30365, C2 =>
                           n29540, A => n27183, ZN => n27170);
   U22821 : OAI22_X1 port map( A1 => n9128, A2 => n30359, B1 => n9896, B2 => 
                           n30353, ZN => n27183);
   U22822 : AOI221_X1 port map( B1 => n30371, B2 => n29733, C1 => n30365, C2 =>
                           n29541, A => n27157, ZN => n27144);
   U22823 : OAI22_X1 port map( A1 => n9123, A2 => n30359, B1 => n9891, B2 => 
                           n30353, ZN => n27157);
   U22824 : AOI221_X1 port map( B1 => n30371, B2 => n29734, C1 => n30365, C2 =>
                           n29542, A => n27131, ZN => n27118);
   U22825 : OAI22_X1 port map( A1 => n9118, A2 => n30359, B1 => n9886, B2 => 
                           n30353, ZN => n27131);
   U22826 : AOI221_X1 port map( B1 => n30371, B2 => n29735, C1 => n30365, C2 =>
                           n29543, A => n27105, ZN => n27092);
   U22827 : OAI22_X1 port map( A1 => n9113, A2 => n30359, B1 => n9881, B2 => 
                           n30353, ZN => n27105);
   U22828 : AOI221_X1 port map( B1 => n30372, B2 => n29736, C1 => n30366, C2 =>
                           n29544, A => n27079, ZN => n27066);
   U22829 : OAI22_X1 port map( A1 => n9108, A2 => n30360, B1 => n9876, B2 => 
                           n30354, ZN => n27079);
   U22830 : AOI221_X1 port map( B1 => n30372, B2 => n29737, C1 => n30366, C2 =>
                           n29545, A => n27053, ZN => n27040);
   U22831 : OAI22_X1 port map( A1 => n9103, A2 => n30360, B1 => n9871, B2 => 
                           n30354, ZN => n27053);
   U22832 : AOI221_X1 port map( B1 => n30372, B2 => n29738, C1 => n30366, C2 =>
                           n29546, A => n27027, ZN => n27014);
   U22833 : OAI22_X1 port map( A1 => n9098, A2 => n30360, B1 => n9866, B2 => 
                           n30354, ZN => n27027);
   U22834 : AOI221_X1 port map( B1 => n30372, B2 => n29739, C1 => n30366, C2 =>
                           n29547, A => n27001, ZN => n26988);
   U22835 : OAI22_X1 port map( A1 => n9093, A2 => n30360, B1 => n9861, B2 => 
                           n30354, ZN => n27001);
   U22836 : AOI221_X1 port map( B1 => n30372, B2 => n29740, C1 => n30366, C2 =>
                           n29548, A => n26975, ZN => n26962);
   U22837 : OAI22_X1 port map( A1 => n9088, A2 => n30360, B1 => n9856, B2 => 
                           n30354, ZN => n26975);
   U22838 : AOI221_X1 port map( B1 => n30372, B2 => n29741, C1 => n30366, C2 =>
                           n29549, A => n26949, ZN => n26936);
   U22839 : OAI22_X1 port map( A1 => n9083, A2 => n30360, B1 => n9851, B2 => 
                           n30354, ZN => n26949);
   U22840 : AOI221_X1 port map( B1 => n30372, B2 => n29742, C1 => n30366, C2 =>
                           n29550, A => n26923, ZN => n26910);
   U22841 : OAI22_X1 port map( A1 => n9078, A2 => n30360, B1 => n9846, B2 => 
                           n30354, ZN => n26923);
   U22842 : AOI221_X1 port map( B1 => n30372, B2 => n29743, C1 => n30366, C2 =>
                           n29551, A => n26897, ZN => n26884);
   U22843 : OAI22_X1 port map( A1 => n9073, A2 => n30360, B1 => n9841, B2 => 
                           n30354, ZN => n26897);
   U22844 : AOI221_X1 port map( B1 => n30372, B2 => n29744, C1 => n30366, C2 =>
                           n29552, A => n26871, ZN => n26858);
   U22845 : OAI22_X1 port map( A1 => n9068, A2 => n30360, B1 => n9836, B2 => 
                           n30354, ZN => n26871);
   U22846 : AOI221_X1 port map( B1 => n30372, B2 => n29745, C1 => n30366, C2 =>
                           n29553, A => n26845, ZN => n26832);
   U22847 : OAI22_X1 port map( A1 => n9063, A2 => n30360, B1 => n9831, B2 => 
                           n30354, ZN => n26845);
   U22848 : AOI221_X1 port map( B1 => n30372, B2 => n29746, C1 => n30366, C2 =>
                           n29554, A => n26819, ZN => n26806);
   U22849 : OAI22_X1 port map( A1 => n9058, A2 => n30360, B1 => n9826, B2 => 
                           n30354, ZN => n26819);
   U22850 : AOI221_X1 port map( B1 => n30372, B2 => n29747, C1 => n30366, C2 =>
                           n29555, A => n26793, ZN => n26780);
   U22851 : OAI22_X1 port map( A1 => n9053, A2 => n30360, B1 => n9821, B2 => 
                           n30354, ZN => n26793);
   U22852 : AOI221_X1 port map( B1 => n30373, B2 => n29748, C1 => n30367, C2 =>
                           n29556, A => n26767, ZN => n26754);
   U22853 : OAI22_X1 port map( A1 => n9048, A2 => n30361, B1 => n9816, B2 => 
                           n30355, ZN => n26767);
   U22854 : AOI221_X1 port map( B1 => n30373, B2 => n29749, C1 => n30367, C2 =>
                           n29557, A => n26741, ZN => n26728);
   U22855 : OAI22_X1 port map( A1 => n9043, A2 => n30361, B1 => n9811, B2 => 
                           n30355, ZN => n26741);
   U22856 : AOI221_X1 port map( B1 => n30373, B2 => n29750, C1 => n30367, C2 =>
                           n29558, A => n26715, ZN => n26702);
   U22857 : OAI22_X1 port map( A1 => n9038, A2 => n30361, B1 => n9806, B2 => 
                           n30355, ZN => n26715);
   U22858 : AOI221_X1 port map( B1 => n30373, B2 => n29751, C1 => n30367, C2 =>
                           n29559, A => n26689, ZN => n26676);
   U22859 : OAI22_X1 port map( A1 => n9033, A2 => n30361, B1 => n9801, B2 => 
                           n30355, ZN => n26689);
   U22860 : AOI221_X1 port map( B1 => n30373, B2 => n29752, C1 => n30367, C2 =>
                           n29560, A => n26663, ZN => n26650);
   U22861 : OAI22_X1 port map( A1 => n9028, A2 => n30361, B1 => n9796, B2 => 
                           n30355, ZN => n26663);
   U22862 : AOI221_X1 port map( B1 => n30373, B2 => n29753, C1 => n30367, C2 =>
                           n29561, A => n26637, ZN => n26624);
   U22863 : OAI22_X1 port map( A1 => n9023, A2 => n30361, B1 => n9791, B2 => 
                           n30355, ZN => n26637);
   U22864 : AOI221_X1 port map( B1 => n30373, B2 => n29754, C1 => n30367, C2 =>
                           n29562, A => n26611, ZN => n26598);
   U22865 : OAI22_X1 port map( A1 => n9018, A2 => n30361, B1 => n9786, B2 => 
                           n30355, ZN => n26611);
   U22866 : AOI221_X1 port map( B1 => n30373, B2 => n29755, C1 => n30367, C2 =>
                           n29563, A => n26585, ZN => n26572);
   U22867 : OAI22_X1 port map( A1 => n9013, A2 => n30361, B1 => n9781, B2 => 
                           n30355, ZN => n26585);
   U22868 : AOI221_X1 port map( B1 => n30373, B2 => n29756, C1 => n30367, C2 =>
                           n29564, A => n26559, ZN => n26546);
   U22869 : OAI22_X1 port map( A1 => n9008, A2 => n30361, B1 => n9776, B2 => 
                           n30355, ZN => n26559);
   U22870 : AOI221_X1 port map( B1 => n30373, B2 => n29757, C1 => n30367, C2 =>
                           n29565, A => n26533, ZN => n26520);
   U22871 : OAI22_X1 port map( A1 => n9003, A2 => n30361, B1 => n9771, B2 => 
                           n30355, ZN => n26533);
   U22872 : AOI221_X1 port map( B1 => n30373, B2 => n29758, C1 => n30367, C2 =>
                           n29566, A => n26507, ZN => n26494);
   U22873 : OAI22_X1 port map( A1 => n8998, A2 => n30361, B1 => n9766, B2 => 
                           n30355, ZN => n26507);
   U22874 : AOI221_X1 port map( B1 => n30373, B2 => n29759, C1 => n30367, C2 =>
                           n29567, A => n26481, ZN => n26468);
   U22875 : OAI22_X1 port map( A1 => n8993, A2 => n30361, B1 => n9761, B2 => 
                           n30355, ZN => n26481);
   U22876 : AOI221_X1 port map( B1 => n30374, B2 => n29760, C1 => n30368, C2 =>
                           n29568, A => n26455, ZN => n26442);
   U22877 : OAI22_X1 port map( A1 => n8988, A2 => n30362, B1 => n9756, B2 => 
                           n30356, ZN => n26455);
   U22878 : AOI221_X1 port map( B1 => n30374, B2 => n29761, C1 => n30368, C2 =>
                           n29569, A => n26429, ZN => n26416);
   U22879 : OAI22_X1 port map( A1 => n8983, A2 => n30362, B1 => n9751, B2 => 
                           n30356, ZN => n26429);
   U22880 : AOI221_X1 port map( B1 => n30374, B2 => n29762, C1 => n30368, C2 =>
                           n29570, A => n26403, ZN => n26390);
   U22881 : OAI22_X1 port map( A1 => n8978, A2 => n30362, B1 => n9746, B2 => 
                           n30356, ZN => n26403);
   U22882 : AOI221_X1 port map( B1 => n30374, B2 => n29763, C1 => n30368, C2 =>
                           n29571, A => n26375, ZN => n26348);
   U22883 : OAI22_X1 port map( A1 => n8973, A2 => n30362, B1 => n9741, B2 => 
                           n30356, ZN => n26375);
   U22884 : NAND2_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(1), ZN => n25451);
   U22885 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => n26100, ZN => n25302);
   U22886 : NAND2_X1 port map( A1 => ADD_WR(2), A2 => n26101, ZN => n25382);
   U22887 : OAI221_X1 port map( B1 => n31124, B2 => n30555, C1 => n31181, C2 =>
                           n10764, A => n26431, ZN => n5889);
   U22888 : OAI21_X1 port map( B1 => n26432, B2 => n26433, A => n30549, ZN => 
                           n26431);
   U22889 : NAND4_X1 port map( A1 => n26442, A2 => n26443, A3 => n26444, A4 => 
                           n26445, ZN => n26432);
   U22890 : NAND4_X1 port map( A1 => n26434, A2 => n26435, A3 => n26436, A4 => 
                           n26437, ZN => n26433);
   U22891 : OAI221_X1 port map( B1 => n31127, B2 => n30555, C1 => n31181, C2 =>
                           n10763, A => n26405, ZN => n5891);
   U22892 : OAI21_X1 port map( B1 => n26406, B2 => n26407, A => n30549, ZN => 
                           n26405);
   U22893 : NAND4_X1 port map( A1 => n26416, A2 => n26417, A3 => n26418, A4 => 
                           n26419, ZN => n26406);
   U22894 : NAND4_X1 port map( A1 => n26408, A2 => n26409, A3 => n26410, A4 => 
                           n26411, ZN => n26407);
   U22895 : OAI221_X1 port map( B1 => n31130, B2 => n30555, C1 => n31181, C2 =>
                           n10762, A => n26379, ZN => n5893);
   U22896 : OAI21_X1 port map( B1 => n26380, B2 => n26381, A => n30549, ZN => 
                           n26379);
   U22897 : NAND4_X1 port map( A1 => n26390, A2 => n26391, A3 => n26392, A4 => 
                           n26393, ZN => n26380);
   U22898 : NAND4_X1 port map( A1 => n26382, A2 => n26383, A3 => n26384, A4 => 
                           n26385, ZN => n26381);
   U22899 : AOI221_X1 port map( B1 => n30495, B2 => n22012, C1 => n30489, C2 =>
                           n9306, A => n26440, ZN => n26435);
   U22900 : OAI22_X1 port map( A1 => n25741, A2 => n30483, B1 => n25675, B2 => 
                           n30477, ZN => n26440);
   U22901 : AOI221_X1 port map( B1 => n30446, B2 => n21919, C1 => n30440, C2 =>
                           n9308, A => n26446, ZN => n26445);
   U22902 : OAI22_X1 port map( A1 => n26028, A2 => n30434, B1 => n25962, B2 => 
                           n30428, ZN => n26446);
   U22903 : AOI221_X1 port map( B1 => n30495, B2 => n22013, C1 => n30489, C2 =>
                           n9301, A => n26414, ZN => n26409);
   U22904 : OAI22_X1 port map( A1 => n25740, A2 => n30483, B1 => n25674, B2 => 
                           n30477, ZN => n26414);
   U22905 : AOI221_X1 port map( B1 => n30446, B2 => n21920, C1 => n30440, C2 =>
                           n9303, A => n26420, ZN => n26419);
   U22906 : OAI22_X1 port map( A1 => n26027, A2 => n30434, B1 => n25961, B2 => 
                           n30428, ZN => n26420);
   U22907 : AOI221_X1 port map( B1 => n30495, B2 => n22014, C1 => n30489, C2 =>
                           n9296, A => n26388, ZN => n26383);
   U22908 : OAI22_X1 port map( A1 => n25739, A2 => n30483, B1 => n25673, B2 => 
                           n30477, ZN => n26388);
   U22909 : AOI221_X1 port map( B1 => n30446, B2 => n21921, C1 => n30440, C2 =>
                           n9298, A => n26394, ZN => n26393);
   U22910 : OAI22_X1 port map( A1 => n26026, A2 => n30434, B1 => n25960, B2 => 
                           n30428, ZN => n26394);
   U22911 : AOI221_X1 port map( B1 => n30495, B2 => n22015, C1 => n30489, C2 =>
                           n9291, A => n26340, ZN => n26325);
   U22912 : OAI22_X1 port map( A1 => n25737, A2 => n30483, B1 => n25671, B2 => 
                           n30477, ZN => n26340);
   U22913 : AOI221_X1 port map( B1 => n30446, B2 => n21922, C1 => n30440, C2 =>
                           n9293, A => n26354, ZN => n26351);
   U22914 : OAI22_X1 port map( A1 => n26024, A2 => n30434, B1 => n25958, B2 => 
                           n30428, ZN => n26354);
   U22915 : OAI221_X1 port map( B1 => n30944, B2 => n30345, C1 => n31180, C2 =>
                           n10888, A => n29272, ZN => n5642);
   U22916 : OAI21_X1 port map( B1 => n29273, B2 => n29274, A => n30339, ZN => 
                           n29272);
   U22917 : NAND4_X1 port map( A1 => n29276, A2 => n29277, A3 => n29278, A4 => 
                           n29279, ZN => n29274);
   U22918 : NAND4_X1 port map( A1 => n29294, A2 => n29295, A3 => n29296, A4 => 
                           n29297, ZN => n29273);
   U22919 : OAI221_X1 port map( B1 => n30947, B2 => n30345, C1 => n31179, C2 =>
                           n10887, A => n29253, ZN => n5644);
   U22920 : OAI21_X1 port map( B1 => n29254, B2 => n29255, A => n30339, ZN => 
                           n29253);
   U22921 : NAND4_X1 port map( A1 => n29256, A2 => n29257, A3 => n29258, A4 => 
                           n29259, ZN => n29255);
   U22922 : NAND4_X1 port map( A1 => n29264, A2 => n29265, A3 => n29266, A4 => 
                           n29267, ZN => n29254);
   U22923 : OAI221_X1 port map( B1 => n30950, B2 => n30345, C1 => n31179, C2 =>
                           n10886, A => n29234, ZN => n5646);
   U22924 : OAI21_X1 port map( B1 => n29235, B2 => n29236, A => n30339, ZN => 
                           n29234);
   U22925 : NAND4_X1 port map( A1 => n29237, A2 => n29238, A3 => n29239, A4 => 
                           n29240, ZN => n29236);
   U22926 : NAND4_X1 port map( A1 => n29245, A2 => n29246, A3 => n29247, A4 => 
                           n29248, ZN => n29235);
   U22927 : OAI221_X1 port map( B1 => n30953, B2 => n30345, C1 => n31179, C2 =>
                           n10885, A => n29215, ZN => n5648);
   U22928 : OAI21_X1 port map( B1 => n29216, B2 => n29217, A => n30339, ZN => 
                           n29215);
   U22929 : NAND4_X1 port map( A1 => n29218, A2 => n29219, A3 => n29220, A4 => 
                           n29221, ZN => n29217);
   U22930 : NAND4_X1 port map( A1 => n29226, A2 => n29227, A3 => n29228, A4 => 
                           n29229, ZN => n29216);
   U22931 : OAI221_X1 port map( B1 => n30956, B2 => n30345, C1 => n31179, C2 =>
                           n10884, A => n29196, ZN => n5650);
   U22932 : OAI21_X1 port map( B1 => n29197, B2 => n29198, A => n30339, ZN => 
                           n29196);
   U22933 : NAND4_X1 port map( A1 => n29199, A2 => n29200, A3 => n29201, A4 => 
                           n29202, ZN => n29198);
   U22934 : NAND4_X1 port map( A1 => n29207, A2 => n29208, A3 => n29209, A4 => 
                           n29210, ZN => n29197);
   U22935 : OAI221_X1 port map( B1 => n30959, B2 => n30345, C1 => n31179, C2 =>
                           n10883, A => n29177, ZN => n5652);
   U22936 : OAI21_X1 port map( B1 => n29178, B2 => n29179, A => n30339, ZN => 
                           n29177);
   U22937 : NAND4_X1 port map( A1 => n29180, A2 => n29181, A3 => n29182, A4 => 
                           n29183, ZN => n29179);
   U22938 : NAND4_X1 port map( A1 => n29188, A2 => n29189, A3 => n29190, A4 => 
                           n29191, ZN => n29178);
   U22939 : OAI221_X1 port map( B1 => n30962, B2 => n30345, C1 => n31179, C2 =>
                           n10882, A => n29158, ZN => n5654);
   U22940 : OAI21_X1 port map( B1 => n29159, B2 => n29160, A => n30339, ZN => 
                           n29158);
   U22941 : NAND4_X1 port map( A1 => n29161, A2 => n29162, A3 => n29163, A4 => 
                           n29164, ZN => n29160);
   U22942 : NAND4_X1 port map( A1 => n29169, A2 => n29170, A3 => n29171, A4 => 
                           n29172, ZN => n29159);
   U22943 : OAI221_X1 port map( B1 => n30965, B2 => n30345, C1 => n31179, C2 =>
                           n10881, A => n29139, ZN => n5656);
   U22944 : OAI21_X1 port map( B1 => n29140, B2 => n29141, A => n30339, ZN => 
                           n29139);
   U22945 : NAND4_X1 port map( A1 => n29142, A2 => n29143, A3 => n29144, A4 => 
                           n29145, ZN => n29141);
   U22946 : NAND4_X1 port map( A1 => n29150, A2 => n29151, A3 => n29152, A4 => 
                           n29153, ZN => n29140);
   U22947 : OAI221_X1 port map( B1 => n30968, B2 => n30345, C1 => n31179, C2 =>
                           n10880, A => n29120, ZN => n5658);
   U22948 : OAI21_X1 port map( B1 => n29121, B2 => n29122, A => n30339, ZN => 
                           n29120);
   U22949 : NAND4_X1 port map( A1 => n29123, A2 => n29124, A3 => n29125, A4 => 
                           n29126, ZN => n29122);
   U22950 : NAND4_X1 port map( A1 => n29131, A2 => n29132, A3 => n29133, A4 => 
                           n29134, ZN => n29121);
   U22951 : OAI221_X1 port map( B1 => n30971, B2 => n30345, C1 => n31179, C2 =>
                           n10879, A => n29101, ZN => n5660);
   U22952 : OAI21_X1 port map( B1 => n29102, B2 => n29103, A => n30339, ZN => 
                           n29101);
   U22953 : NAND4_X1 port map( A1 => n29104, A2 => n29105, A3 => n29106, A4 => 
                           n29107, ZN => n29103);
   U22954 : NAND4_X1 port map( A1 => n29112, A2 => n29113, A3 => n29114, A4 => 
                           n29115, ZN => n29102);
   U22955 : OAI221_X1 port map( B1 => n30974, B2 => n30345, C1 => n31179, C2 =>
                           n10878, A => n29082, ZN => n5662);
   U22956 : OAI21_X1 port map( B1 => n29083, B2 => n29084, A => n30339, ZN => 
                           n29082);
   U22957 : NAND4_X1 port map( A1 => n29085, A2 => n29086, A3 => n29087, A4 => 
                           n29088, ZN => n29084);
   U22958 : NAND4_X1 port map( A1 => n29093, A2 => n29094, A3 => n29095, A4 => 
                           n29096, ZN => n29083);
   U22959 : OAI221_X1 port map( B1 => n30977, B2 => n30345, C1 => n31179, C2 =>
                           n10877, A => n29063, ZN => n5664);
   U22960 : OAI21_X1 port map( B1 => n29064, B2 => n29065, A => n30339, ZN => 
                           n29063);
   U22961 : NAND4_X1 port map( A1 => n29066, A2 => n29067, A3 => n29068, A4 => 
                           n29069, ZN => n29065);
   U22962 : NAND4_X1 port map( A1 => n29074, A2 => n29075, A3 => n29076, A4 => 
                           n29077, ZN => n29064);
   U22963 : OAI221_X1 port map( B1 => n30980, B2 => n30346, C1 => n31179, C2 =>
                           n10876, A => n29044, ZN => n5666);
   U22964 : OAI21_X1 port map( B1 => n29045, B2 => n29046, A => n30340, ZN => 
                           n29044);
   U22965 : NAND4_X1 port map( A1 => n29047, A2 => n29048, A3 => n29049, A4 => 
                           n29050, ZN => n29046);
   U22966 : NAND4_X1 port map( A1 => n29055, A2 => n29056, A3 => n29057, A4 => 
                           n29058, ZN => n29045);
   U22967 : OAI221_X1 port map( B1 => n30983, B2 => n30346, C1 => n31180, C2 =>
                           n10875, A => n29025, ZN => n5668);
   U22968 : OAI21_X1 port map( B1 => n29026, B2 => n29027, A => n30340, ZN => 
                           n29025);
   U22969 : NAND4_X1 port map( A1 => n29028, A2 => n29029, A3 => n29030, A4 => 
                           n29031, ZN => n29027);
   U22970 : NAND4_X1 port map( A1 => n29036, A2 => n29037, A3 => n29038, A4 => 
                           n29039, ZN => n29026);
   U22971 : OAI221_X1 port map( B1 => n30986, B2 => n30346, C1 => n31178, C2 =>
                           n10874, A => n29006, ZN => n5670);
   U22972 : OAI21_X1 port map( B1 => n29007, B2 => n29008, A => n30340, ZN => 
                           n29006);
   U22973 : NAND4_X1 port map( A1 => n29009, A2 => n29010, A3 => n29011, A4 => 
                           n29012, ZN => n29008);
   U22974 : NAND4_X1 port map( A1 => n29017, A2 => n29018, A3 => n29019, A4 => 
                           n29020, ZN => n29007);
   U22975 : OAI221_X1 port map( B1 => n30989, B2 => n30346, C1 => n31178, C2 =>
                           n10873, A => n28987, ZN => n5672);
   U22976 : OAI21_X1 port map( B1 => n28988, B2 => n28989, A => n30340, ZN => 
                           n28987);
   U22977 : NAND4_X1 port map( A1 => n28990, A2 => n28991, A3 => n28992, A4 => 
                           n28993, ZN => n28989);
   U22978 : NAND4_X1 port map( A1 => n28998, A2 => n28999, A3 => n29000, A4 => 
                           n29001, ZN => n28988);
   U22979 : OAI221_X1 port map( B1 => n30992, B2 => n30346, C1 => n31178, C2 =>
                           n10872, A => n28968, ZN => n5674);
   U22980 : OAI21_X1 port map( B1 => n28969, B2 => n28970, A => n30340, ZN => 
                           n28968);
   U22981 : NAND4_X1 port map( A1 => n28971, A2 => n28972, A3 => n28973, A4 => 
                           n28974, ZN => n28970);
   U22982 : NAND4_X1 port map( A1 => n28979, A2 => n28980, A3 => n28981, A4 => 
                           n28982, ZN => n28969);
   U22983 : OAI221_X1 port map( B1 => n30995, B2 => n30346, C1 => n31178, C2 =>
                           n10871, A => n28949, ZN => n5676);
   U22984 : OAI21_X1 port map( B1 => n28950, B2 => n28951, A => n30340, ZN => 
                           n28949);
   U22985 : NAND4_X1 port map( A1 => n28952, A2 => n28953, A3 => n28954, A4 => 
                           n28955, ZN => n28951);
   U22986 : NAND4_X1 port map( A1 => n28960, A2 => n28961, A3 => n28962, A4 => 
                           n28963, ZN => n28950);
   U22987 : OAI221_X1 port map( B1 => n30998, B2 => n30346, C1 => n31178, C2 =>
                           n10870, A => n28930, ZN => n5678);
   U22988 : OAI21_X1 port map( B1 => n28931, B2 => n28932, A => n30340, ZN => 
                           n28930);
   U22989 : NAND4_X1 port map( A1 => n28933, A2 => n28934, A3 => n28935, A4 => 
                           n28936, ZN => n28932);
   U22990 : NAND4_X1 port map( A1 => n28941, A2 => n28942, A3 => n28943, A4 => 
                           n28944, ZN => n28931);
   U22991 : OAI221_X1 port map( B1 => n31001, B2 => n30346, C1 => n31178, C2 =>
                           n10869, A => n28911, ZN => n5680);
   U22992 : OAI21_X1 port map( B1 => n28912, B2 => n28913, A => n30340, ZN => 
                           n28911);
   U22993 : NAND4_X1 port map( A1 => n28914, A2 => n28915, A3 => n28916, A4 => 
                           n28917, ZN => n28913);
   U22994 : NAND4_X1 port map( A1 => n28922, A2 => n28923, A3 => n28924, A4 => 
                           n28925, ZN => n28912);
   U22995 : OAI221_X1 port map( B1 => n31004, B2 => n30346, C1 => n31178, C2 =>
                           n10868, A => n28892, ZN => n5682);
   U22996 : OAI21_X1 port map( B1 => n28893, B2 => n28894, A => n30340, ZN => 
                           n28892);
   U22997 : NAND4_X1 port map( A1 => n28895, A2 => n28896, A3 => n28897, A4 => 
                           n28898, ZN => n28894);
   U22998 : NAND4_X1 port map( A1 => n28903, A2 => n28904, A3 => n28905, A4 => 
                           n28906, ZN => n28893);
   U22999 : OAI221_X1 port map( B1 => n31007, B2 => n30346, C1 => n31178, C2 =>
                           n10867, A => n28873, ZN => n5684);
   U23000 : OAI21_X1 port map( B1 => n28874, B2 => n28875, A => n30340, ZN => 
                           n28873);
   U23001 : NAND4_X1 port map( A1 => n28876, A2 => n28877, A3 => n28878, A4 => 
                           n28879, ZN => n28875);
   U23002 : NAND4_X1 port map( A1 => n28884, A2 => n28885, A3 => n28886, A4 => 
                           n28887, ZN => n28874);
   U23003 : OAI221_X1 port map( B1 => n31010, B2 => n30346, C1 => n31178, C2 =>
                           n10866, A => n28854, ZN => n5686);
   U23004 : OAI21_X1 port map( B1 => n28855, B2 => n28856, A => n30340, ZN => 
                           n28854);
   U23005 : NAND4_X1 port map( A1 => n28857, A2 => n28858, A3 => n28859, A4 => 
                           n28860, ZN => n28856);
   U23006 : NAND4_X1 port map( A1 => n28865, A2 => n28866, A3 => n28867, A4 => 
                           n28868, ZN => n28855);
   U23007 : OAI221_X1 port map( B1 => n31013, B2 => n30346, C1 => n31178, C2 =>
                           n10865, A => n28835, ZN => n5688);
   U23008 : OAI21_X1 port map( B1 => n28836, B2 => n28837, A => n30340, ZN => 
                           n28835);
   U23009 : NAND4_X1 port map( A1 => n28838, A2 => n28839, A3 => n28840, A4 => 
                           n28841, ZN => n28837);
   U23010 : NAND4_X1 port map( A1 => n28846, A2 => n28847, A3 => n28848, A4 => 
                           n28849, ZN => n28836);
   U23011 : OAI221_X1 port map( B1 => n31016, B2 => n30347, C1 => n31178, C2 =>
                           n10864, A => n28816, ZN => n5690);
   U23012 : OAI21_X1 port map( B1 => n28817, B2 => n28818, A => n30341, ZN => 
                           n28816);
   U23013 : NAND4_X1 port map( A1 => n28819, A2 => n28820, A3 => n28821, A4 => 
                           n28822, ZN => n28818);
   U23014 : NAND4_X1 port map( A1 => n28827, A2 => n28828, A3 => n28829, A4 => 
                           n28830, ZN => n28817);
   U23015 : OAI221_X1 port map( B1 => n31019, B2 => n30347, C1 => n31178, C2 =>
                           n10863, A => n28797, ZN => n5692);
   U23016 : OAI21_X1 port map( B1 => n28798, B2 => n28799, A => n30341, ZN => 
                           n28797);
   U23017 : NAND4_X1 port map( A1 => n28800, A2 => n28801, A3 => n28802, A4 => 
                           n28803, ZN => n28799);
   U23018 : NAND4_X1 port map( A1 => n28808, A2 => n28809, A3 => n28810, A4 => 
                           n28811, ZN => n28798);
   U23019 : OAI221_X1 port map( B1 => n31022, B2 => n30347, C1 => n31177, C2 =>
                           n10862, A => n28778, ZN => n5694);
   U23020 : OAI21_X1 port map( B1 => n28779, B2 => n28780, A => n30341, ZN => 
                           n28778);
   U23021 : NAND4_X1 port map( A1 => n28781, A2 => n28782, A3 => n28783, A4 => 
                           n28784, ZN => n28780);
   U23022 : NAND4_X1 port map( A1 => n28789, A2 => n28790, A3 => n28791, A4 => 
                           n28792, ZN => n28779);
   U23023 : OAI221_X1 port map( B1 => n31025, B2 => n30347, C1 => n31177, C2 =>
                           n10861, A => n28759, ZN => n5696);
   U23024 : OAI21_X1 port map( B1 => n28760, B2 => n28761, A => n30341, ZN => 
                           n28759);
   U23025 : NAND4_X1 port map( A1 => n28762, A2 => n28763, A3 => n28764, A4 => 
                           n28765, ZN => n28761);
   U23026 : NAND4_X1 port map( A1 => n28770, A2 => n28771, A3 => n28772, A4 => 
                           n28773, ZN => n28760);
   U23027 : OAI221_X1 port map( B1 => n31028, B2 => n30347, C1 => n31177, C2 =>
                           n10860, A => n28740, ZN => n5698);
   U23028 : OAI21_X1 port map( B1 => n28741, B2 => n28742, A => n30341, ZN => 
                           n28740);
   U23029 : NAND4_X1 port map( A1 => n28743, A2 => n28744, A3 => n28745, A4 => 
                           n28746, ZN => n28742);
   U23030 : NAND4_X1 port map( A1 => n28751, A2 => n28752, A3 => n28753, A4 => 
                           n28754, ZN => n28741);
   U23031 : OAI221_X1 port map( B1 => n31031, B2 => n30347, C1 => n31177, C2 =>
                           n10859, A => n28721, ZN => n5700);
   U23032 : OAI21_X1 port map( B1 => n28722, B2 => n28723, A => n30341, ZN => 
                           n28721);
   U23033 : NAND4_X1 port map( A1 => n28724, A2 => n28725, A3 => n28726, A4 => 
                           n28727, ZN => n28723);
   U23034 : NAND4_X1 port map( A1 => n28732, A2 => n28733, A3 => n28734, A4 => 
                           n28735, ZN => n28722);
   U23035 : OAI221_X1 port map( B1 => n31034, B2 => n30347, C1 => n31177, C2 =>
                           n10858, A => n28702, ZN => n5702);
   U23036 : OAI21_X1 port map( B1 => n28703, B2 => n28704, A => n30341, ZN => 
                           n28702);
   U23037 : NAND4_X1 port map( A1 => n28705, A2 => n28706, A3 => n28707, A4 => 
                           n28708, ZN => n28704);
   U23038 : NAND4_X1 port map( A1 => n28713, A2 => n28714, A3 => n28715, A4 => 
                           n28716, ZN => n28703);
   U23039 : OAI221_X1 port map( B1 => n31037, B2 => n30347, C1 => n31177, C2 =>
                           n10857, A => n28683, ZN => n5704);
   U23040 : OAI21_X1 port map( B1 => n28684, B2 => n28685, A => n30341, ZN => 
                           n28683);
   U23041 : NAND4_X1 port map( A1 => n28686, A2 => n28687, A3 => n28688, A4 => 
                           n28689, ZN => n28685);
   U23042 : NAND4_X1 port map( A1 => n28694, A2 => n28695, A3 => n28696, A4 => 
                           n28697, ZN => n28684);
   U23043 : OAI221_X1 port map( B1 => n31040, B2 => n30347, C1 => n31177, C2 =>
                           n10856, A => n28664, ZN => n5706);
   U23044 : OAI21_X1 port map( B1 => n28665, B2 => n28666, A => n30341, ZN => 
                           n28664);
   U23045 : NAND4_X1 port map( A1 => n28667, A2 => n28668, A3 => n28669, A4 => 
                           n28670, ZN => n28666);
   U23046 : NAND4_X1 port map( A1 => n28675, A2 => n28676, A3 => n28677, A4 => 
                           n28678, ZN => n28665);
   U23047 : OAI221_X1 port map( B1 => n31043, B2 => n30347, C1 => n31177, C2 =>
                           n10855, A => n28645, ZN => n5708);
   U23048 : OAI21_X1 port map( B1 => n28646, B2 => n28647, A => n30341, ZN => 
                           n28645);
   U23049 : NAND4_X1 port map( A1 => n28648, A2 => n28649, A3 => n28650, A4 => 
                           n28651, ZN => n28647);
   U23050 : NAND4_X1 port map( A1 => n28656, A2 => n28657, A3 => n28658, A4 => 
                           n28659, ZN => n28646);
   U23051 : OAI221_X1 port map( B1 => n31046, B2 => n30347, C1 => n31177, C2 =>
                           n10854, A => n28626, ZN => n5710);
   U23052 : OAI21_X1 port map( B1 => n28627, B2 => n28628, A => n30341, ZN => 
                           n28626);
   U23053 : NAND4_X1 port map( A1 => n28629, A2 => n28630, A3 => n28631, A4 => 
                           n28632, ZN => n28628);
   U23054 : NAND4_X1 port map( A1 => n28637, A2 => n28638, A3 => n28639, A4 => 
                           n28640, ZN => n28627);
   U23055 : OAI221_X1 port map( B1 => n31049, B2 => n30347, C1 => n31177, C2 =>
                           n10853, A => n28607, ZN => n5712);
   U23056 : OAI21_X1 port map( B1 => n28608, B2 => n28609, A => n30341, ZN => 
                           n28607);
   U23057 : NAND4_X1 port map( A1 => n28610, A2 => n28611, A3 => n28612, A4 => 
                           n28613, ZN => n28609);
   U23058 : NAND4_X1 port map( A1 => n28618, A2 => n28619, A3 => n28620, A4 => 
                           n28621, ZN => n28608);
   U23059 : OAI221_X1 port map( B1 => n31052, B2 => n30348, C1 => n31177, C2 =>
                           n10852, A => n28588, ZN => n5714);
   U23060 : OAI21_X1 port map( B1 => n28589, B2 => n28590, A => n30342, ZN => 
                           n28588);
   U23061 : NAND4_X1 port map( A1 => n28591, A2 => n28592, A3 => n28593, A4 => 
                           n28594, ZN => n28590);
   U23062 : NAND4_X1 port map( A1 => n28599, A2 => n28600, A3 => n28601, A4 => 
                           n28602, ZN => n28589);
   U23063 : OAI221_X1 port map( B1 => n31055, B2 => n30348, C1 => n31178, C2 =>
                           n10851, A => n28569, ZN => n5716);
   U23064 : OAI21_X1 port map( B1 => n28570, B2 => n28571, A => n30342, ZN => 
                           n28569);
   U23065 : NAND4_X1 port map( A1 => n28572, A2 => n28573, A3 => n28574, A4 => 
                           n28575, ZN => n28571);
   U23066 : NAND4_X1 port map( A1 => n28580, A2 => n28581, A3 => n28582, A4 => 
                           n28583, ZN => n28570);
   U23067 : OAI221_X1 port map( B1 => n31058, B2 => n30348, C1 => n31179, C2 =>
                           n10850, A => n28550, ZN => n5718);
   U23068 : OAI21_X1 port map( B1 => n28551, B2 => n28552, A => n30342, ZN => 
                           n28550);
   U23069 : NAND4_X1 port map( A1 => n28553, A2 => n28554, A3 => n28555, A4 => 
                           n28556, ZN => n28552);
   U23070 : NAND4_X1 port map( A1 => n28561, A2 => n28562, A3 => n28563, A4 => 
                           n28564, ZN => n28551);
   U23071 : OAI221_X1 port map( B1 => n31061, B2 => n30348, C1 => n31180, C2 =>
                           n10849, A => n28531, ZN => n5720);
   U23072 : OAI21_X1 port map( B1 => n28532, B2 => n28533, A => n30342, ZN => 
                           n28531);
   U23073 : NAND4_X1 port map( A1 => n28534, A2 => n28535, A3 => n28536, A4 => 
                           n28537, ZN => n28533);
   U23074 : NAND4_X1 port map( A1 => n28542, A2 => n28543, A3 => n28544, A4 => 
                           n28545, ZN => n28532);
   U23075 : OAI221_X1 port map( B1 => n31064, B2 => n30348, C1 => n31180, C2 =>
                           n10848, A => n28512, ZN => n5722);
   U23076 : OAI21_X1 port map( B1 => n28513, B2 => n28514, A => n30342, ZN => 
                           n28512);
   U23077 : NAND4_X1 port map( A1 => n28515, A2 => n28516, A3 => n28517, A4 => 
                           n28518, ZN => n28514);
   U23078 : NAND4_X1 port map( A1 => n28523, A2 => n28524, A3 => n28525, A4 => 
                           n28526, ZN => n28513);
   U23079 : OAI221_X1 port map( B1 => n31067, B2 => n30348, C1 => n31180, C2 =>
                           n10847, A => n28493, ZN => n5724);
   U23080 : OAI21_X1 port map( B1 => n28494, B2 => n28495, A => n30342, ZN => 
                           n28493);
   U23081 : NAND4_X1 port map( A1 => n28496, A2 => n28497, A3 => n28498, A4 => 
                           n28499, ZN => n28495);
   U23082 : NAND4_X1 port map( A1 => n28504, A2 => n28505, A3 => n28506, A4 => 
                           n28507, ZN => n28494);
   U23083 : OAI221_X1 port map( B1 => n31070, B2 => n30348, C1 => n31180, C2 =>
                           n10846, A => n28474, ZN => n5726);
   U23084 : OAI21_X1 port map( B1 => n28475, B2 => n28476, A => n30342, ZN => 
                           n28474);
   U23085 : NAND4_X1 port map( A1 => n28477, A2 => n28478, A3 => n28479, A4 => 
                           n28480, ZN => n28476);
   U23086 : NAND4_X1 port map( A1 => n28485, A2 => n28486, A3 => n28487, A4 => 
                           n28488, ZN => n28475);
   U23087 : OAI221_X1 port map( B1 => n31073, B2 => n30348, C1 => n31180, C2 =>
                           n10845, A => n28455, ZN => n5728);
   U23088 : OAI21_X1 port map( B1 => n28456, B2 => n28457, A => n30342, ZN => 
                           n28455);
   U23089 : NAND4_X1 port map( A1 => n28458, A2 => n28459, A3 => n28460, A4 => 
                           n28461, ZN => n28457);
   U23090 : NAND4_X1 port map( A1 => n28466, A2 => n28467, A3 => n28468, A4 => 
                           n28469, ZN => n28456);
   U23091 : OAI221_X1 port map( B1 => n31076, B2 => n30348, C1 => n31180, C2 =>
                           n10844, A => n28436, ZN => n5730);
   U23092 : OAI21_X1 port map( B1 => n28437, B2 => n28438, A => n30342, ZN => 
                           n28436);
   U23093 : NAND4_X1 port map( A1 => n28439, A2 => n28440, A3 => n28441, A4 => 
                           n28442, ZN => n28438);
   U23094 : NAND4_X1 port map( A1 => n28447, A2 => n28448, A3 => n28449, A4 => 
                           n28450, ZN => n28437);
   U23095 : OAI221_X1 port map( B1 => n31079, B2 => n30348, C1 => n31180, C2 =>
                           n10843, A => n28417, ZN => n5732);
   U23096 : OAI21_X1 port map( B1 => n28418, B2 => n28419, A => n30342, ZN => 
                           n28417);
   U23097 : NAND4_X1 port map( A1 => n28420, A2 => n28421, A3 => n28422, A4 => 
                           n28423, ZN => n28419);
   U23098 : NAND4_X1 port map( A1 => n28428, A2 => n28429, A3 => n28430, A4 => 
                           n28431, ZN => n28418);
   U23099 : OAI221_X1 port map( B1 => n31082, B2 => n30348, C1 => n31180, C2 =>
                           n10842, A => n28398, ZN => n5734);
   U23100 : OAI21_X1 port map( B1 => n28399, B2 => n28400, A => n30342, ZN => 
                           n28398);
   U23101 : NAND4_X1 port map( A1 => n28401, A2 => n28402, A3 => n28403, A4 => 
                           n28404, ZN => n28400);
   U23102 : NAND4_X1 port map( A1 => n28409, A2 => n28410, A3 => n28411, A4 => 
                           n28412, ZN => n28399);
   U23103 : OAI221_X1 port map( B1 => n31085, B2 => n30348, C1 => n31180, C2 =>
                           n10841, A => n28379, ZN => n5736);
   U23104 : OAI21_X1 port map( B1 => n28380, B2 => n28381, A => n30342, ZN => 
                           n28379);
   U23105 : NAND4_X1 port map( A1 => n28382, A2 => n28383, A3 => n28384, A4 => 
                           n28385, ZN => n28381);
   U23106 : NAND4_X1 port map( A1 => n28390, A2 => n28391, A3 => n28392, A4 => 
                           n28393, ZN => n28380);
   U23107 : OAI221_X1 port map( B1 => n31088, B2 => n30349, C1 => n31186, C2 =>
                           n10840, A => n28360, ZN => n5738);
   U23108 : OAI21_X1 port map( B1 => n28361, B2 => n28362, A => n30343, ZN => 
                           n28360);
   U23109 : NAND4_X1 port map( A1 => n28363, A2 => n28364, A3 => n28365, A4 => 
                           n28366, ZN => n28362);
   U23110 : NAND4_X1 port map( A1 => n28371, A2 => n28372, A3 => n28373, A4 => 
                           n28374, ZN => n28361);
   U23111 : OAI221_X1 port map( B1 => n31091, B2 => n30349, C1 => n31186, C2 =>
                           n10839, A => n28341, ZN => n5740);
   U23112 : OAI21_X1 port map( B1 => n28342, B2 => n28343, A => n30343, ZN => 
                           n28341);
   U23113 : NAND4_X1 port map( A1 => n28344, A2 => n28345, A3 => n28346, A4 => 
                           n28347, ZN => n28343);
   U23114 : NAND4_X1 port map( A1 => n28352, A2 => n28353, A3 => n28354, A4 => 
                           n28355, ZN => n28342);
   U23115 : OAI221_X1 port map( B1 => n31094, B2 => n30349, C1 => n31186, C2 =>
                           n10838, A => n28322, ZN => n5742);
   U23116 : OAI21_X1 port map( B1 => n28323, B2 => n28324, A => n30343, ZN => 
                           n28322);
   U23117 : NAND4_X1 port map( A1 => n28325, A2 => n28326, A3 => n28327, A4 => 
                           n28328, ZN => n28324);
   U23118 : NAND4_X1 port map( A1 => n28333, A2 => n28334, A3 => n28335, A4 => 
                           n28336, ZN => n28323);
   U23119 : OAI221_X1 port map( B1 => n31097, B2 => n30349, C1 => n31186, C2 =>
                           n10837, A => n28303, ZN => n5744);
   U23120 : OAI21_X1 port map( B1 => n28304, B2 => n28305, A => n30343, ZN => 
                           n28303);
   U23121 : NAND4_X1 port map( A1 => n28306, A2 => n28307, A3 => n28308, A4 => 
                           n28309, ZN => n28305);
   U23122 : NAND4_X1 port map( A1 => n28314, A2 => n28315, A3 => n28316, A4 => 
                           n28317, ZN => n28304);
   U23123 : OAI221_X1 port map( B1 => n31100, B2 => n30349, C1 => n31186, C2 =>
                           n10836, A => n28284, ZN => n5746);
   U23124 : OAI21_X1 port map( B1 => n28285, B2 => n28286, A => n30343, ZN => 
                           n28284);
   U23125 : NAND4_X1 port map( A1 => n28287, A2 => n28288, A3 => n28289, A4 => 
                           n28290, ZN => n28286);
   U23126 : NAND4_X1 port map( A1 => n28295, A2 => n28296, A3 => n28297, A4 => 
                           n28298, ZN => n28285);
   U23127 : OAI221_X1 port map( B1 => n31103, B2 => n30349, C1 => n31180, C2 =>
                           n10835, A => n28265, ZN => n5748);
   U23128 : OAI21_X1 port map( B1 => n28266, B2 => n28267, A => n30343, ZN => 
                           n28265);
   U23129 : NAND4_X1 port map( A1 => n28268, A2 => n28269, A3 => n28270, A4 => 
                           n28271, ZN => n28267);
   U23130 : NAND4_X1 port map( A1 => n28276, A2 => n28277, A3 => n28278, A4 => 
                           n28279, ZN => n28266);
   U23131 : OAI221_X1 port map( B1 => n31106, B2 => n30349, C1 => n31186, C2 =>
                           n10834, A => n28246, ZN => n5750);
   U23132 : OAI21_X1 port map( B1 => n28247, B2 => n28248, A => n30343, ZN => 
                           n28246);
   U23133 : NAND4_X1 port map( A1 => n28249, A2 => n28250, A3 => n28251, A4 => 
                           n28252, ZN => n28248);
   U23134 : NAND4_X1 port map( A1 => n28257, A2 => n28258, A3 => n28259, A4 => 
                           n28260, ZN => n28247);
   U23135 : OAI221_X1 port map( B1 => n31109, B2 => n30349, C1 => n31186, C2 =>
                           n10833, A => n28227, ZN => n5752);
   U23136 : OAI21_X1 port map( B1 => n28228, B2 => n28229, A => n30343, ZN => 
                           n28227);
   U23137 : NAND4_X1 port map( A1 => n28230, A2 => n28231, A3 => n28232, A4 => 
                           n28233, ZN => n28229);
   U23138 : NAND4_X1 port map( A1 => n28238, A2 => n28239, A3 => n28240, A4 => 
                           n28241, ZN => n28228);
   U23139 : OAI221_X1 port map( B1 => n31112, B2 => n30349, C1 => n31186, C2 =>
                           n10832, A => n28208, ZN => n5754);
   U23140 : OAI21_X1 port map( B1 => n28209, B2 => n28210, A => n30343, ZN => 
                           n28208);
   U23141 : NAND4_X1 port map( A1 => n28211, A2 => n28212, A3 => n28213, A4 => 
                           n28214, ZN => n28210);
   U23142 : NAND4_X1 port map( A1 => n28219, A2 => n28220, A3 => n28221, A4 => 
                           n28222, ZN => n28209);
   U23143 : OAI221_X1 port map( B1 => n31115, B2 => n30349, C1 => n31186, C2 =>
                           n10831, A => n28189, ZN => n5756);
   U23144 : OAI21_X1 port map( B1 => n28190, B2 => n28191, A => n30343, ZN => 
                           n28189);
   U23145 : NAND4_X1 port map( A1 => n28192, A2 => n28193, A3 => n28194, A4 => 
                           n28195, ZN => n28191);
   U23146 : NAND4_X1 port map( A1 => n28200, A2 => n28201, A3 => n28202, A4 => 
                           n28203, ZN => n28190);
   U23147 : OAI221_X1 port map( B1 => n31118, B2 => n30349, C1 => n31186, C2 =>
                           n10830, A => n28170, ZN => n5758);
   U23148 : OAI21_X1 port map( B1 => n28171, B2 => n28172, A => n30343, ZN => 
                           n28170);
   U23149 : NAND4_X1 port map( A1 => n28173, A2 => n28174, A3 => n28175, A4 => 
                           n28176, ZN => n28172);
   U23150 : NAND4_X1 port map( A1 => n28181, A2 => n28182, A3 => n28183, A4 => 
                           n28184, ZN => n28171);
   U23151 : OAI221_X1 port map( B1 => n31121, B2 => n30349, C1 => n31186, C2 =>
                           n10829, A => n28151, ZN => n5760);
   U23152 : OAI21_X1 port map( B1 => n28152, B2 => n28153, A => n30343, ZN => 
                           n28151);
   U23153 : NAND4_X1 port map( A1 => n28154, A2 => n28155, A3 => n28156, A4 => 
                           n28157, ZN => n28153);
   U23154 : NAND4_X1 port map( A1 => n28162, A2 => n28163, A3 => n28164, A4 => 
                           n28165, ZN => n28152);
   U23155 : AOI221_X1 port map( B1 => n30285, B2 => n22179, C1 => n30279, C2 =>
                           n9736, A => n29289, ZN => n29277);
   U23156 : OAI22_X1 port map( A1 => n9672, A2 => n30273, B1 => n17836, B2 => 
                           n30267, ZN => n29289);
   U23157 : AOI221_X1 port map( B1 => n30285, B2 => n22180, C1 => n30279, C2 =>
                           n9735, A => n29262, ZN => n29257);
   U23158 : OAI22_X1 port map( A1 => n9671, A2 => n30273, B1 => n17835, B2 => 
                           n30267, ZN => n29262);
   U23159 : AOI221_X1 port map( B1 => n30285, B2 => n22181, C1 => n30279, C2 =>
                           n9734, A => n29243, ZN => n29238);
   U23160 : OAI22_X1 port map( A1 => n9670, A2 => n30273, B1 => n17834, B2 => 
                           n30267, ZN => n29243);
   U23161 : AOI221_X1 port map( B1 => n30285, B2 => n22182, C1 => n30279, C2 =>
                           n9733, A => n29224, ZN => n29219);
   U23162 : OAI22_X1 port map( A1 => n9669, A2 => n30273, B1 => n17833, B2 => 
                           n30267, ZN => n29224);
   U23163 : AOI221_X1 port map( B1 => n30285, B2 => n22183, C1 => n30279, C2 =>
                           n9732, A => n29205, ZN => n29200);
   U23164 : OAI22_X1 port map( A1 => n9668, A2 => n30273, B1 => n17832, B2 => 
                           n30267, ZN => n29205);
   U23165 : AOI221_X1 port map( B1 => n30285, B2 => n22184, C1 => n30279, C2 =>
                           n9731, A => n29186, ZN => n29181);
   U23166 : OAI22_X1 port map( A1 => n9667, A2 => n30273, B1 => n17831, B2 => 
                           n30267, ZN => n29186);
   U23167 : AOI221_X1 port map( B1 => n30285, B2 => n22185, C1 => n30279, C2 =>
                           n9730, A => n29167, ZN => n29162);
   U23168 : OAI22_X1 port map( A1 => n9666, A2 => n30273, B1 => n17830, B2 => 
                           n30267, ZN => n29167);
   U23169 : AOI221_X1 port map( B1 => n30285, B2 => n22186, C1 => n30279, C2 =>
                           n9729, A => n29148, ZN => n29143);
   U23170 : OAI22_X1 port map( A1 => n9665, A2 => n30273, B1 => n17829, B2 => 
                           n30267, ZN => n29148);
   U23171 : AOI221_X1 port map( B1 => n30285, B2 => n22187, C1 => n30279, C2 =>
                           n9728, A => n29129, ZN => n29124);
   U23172 : OAI22_X1 port map( A1 => n9664, A2 => n30273, B1 => n17828, B2 => 
                           n30267, ZN => n29129);
   U23173 : AOI221_X1 port map( B1 => n30285, B2 => n22188, C1 => n30279, C2 =>
                           n9727, A => n29110, ZN => n29105);
   U23174 : OAI22_X1 port map( A1 => n9663, A2 => n30273, B1 => n17827, B2 => 
                           n30267, ZN => n29110);
   U23175 : AOI221_X1 port map( B1 => n30285, B2 => n22189, C1 => n30279, C2 =>
                           n9726, A => n29091, ZN => n29086);
   U23176 : OAI22_X1 port map( A1 => n9662, A2 => n30273, B1 => n17826, B2 => 
                           n30267, ZN => n29091);
   U23177 : AOI221_X1 port map( B1 => n30285, B2 => n22190, C1 => n30279, C2 =>
                           n9725, A => n29072, ZN => n29067);
   U23178 : OAI22_X1 port map( A1 => n9661, A2 => n30273, B1 => n17825, B2 => 
                           n30267, ZN => n29072);
   U23179 : AOI221_X1 port map( B1 => n30286, B2 => n22191, C1 => n30280, C2 =>
                           n9724, A => n29053, ZN => n29048);
   U23180 : OAI22_X1 port map( A1 => n9660, A2 => n30274, B1 => n17824, B2 => 
                           n30268, ZN => n29053);
   U23181 : AOI221_X1 port map( B1 => n30286, B2 => n22192, C1 => n30280, C2 =>
                           n9723, A => n29034, ZN => n29029);
   U23182 : OAI22_X1 port map( A1 => n9659, A2 => n30274, B1 => n17823, B2 => 
                           n30268, ZN => n29034);
   U23183 : AOI221_X1 port map( B1 => n30286, B2 => n22193, C1 => n30280, C2 =>
                           n9722, A => n29015, ZN => n29010);
   U23184 : OAI22_X1 port map( A1 => n9658, A2 => n30274, B1 => n17822, B2 => 
                           n30268, ZN => n29015);
   U23185 : AOI221_X1 port map( B1 => n30286, B2 => n22194, C1 => n30280, C2 =>
                           n9721, A => n28996, ZN => n28991);
   U23186 : OAI22_X1 port map( A1 => n9657, A2 => n30274, B1 => n17821, B2 => 
                           n30268, ZN => n28996);
   U23187 : AOI221_X1 port map( B1 => n30286, B2 => n22195, C1 => n30280, C2 =>
                           n9720, A => n28977, ZN => n28972);
   U23188 : OAI22_X1 port map( A1 => n9656, A2 => n30274, B1 => n17820, B2 => 
                           n30268, ZN => n28977);
   U23189 : AOI221_X1 port map( B1 => n30286, B2 => n22196, C1 => n30280, C2 =>
                           n9719, A => n28958, ZN => n28953);
   U23190 : OAI22_X1 port map( A1 => n9655, A2 => n30274, B1 => n17819, B2 => 
                           n30268, ZN => n28958);
   U23191 : AOI221_X1 port map( B1 => n30286, B2 => n22197, C1 => n30280, C2 =>
                           n9718, A => n28939, ZN => n28934);
   U23192 : OAI22_X1 port map( A1 => n9654, A2 => n30274, B1 => n17818, B2 => 
                           n30268, ZN => n28939);
   U23193 : AOI221_X1 port map( B1 => n30286, B2 => n22198, C1 => n30280, C2 =>
                           n9717, A => n28920, ZN => n28915);
   U23194 : OAI22_X1 port map( A1 => n9653, A2 => n30274, B1 => n17817, B2 => 
                           n30268, ZN => n28920);
   U23195 : AOI221_X1 port map( B1 => n30286, B2 => n22199, C1 => n30280, C2 =>
                           n9716, A => n28901, ZN => n28896);
   U23196 : OAI22_X1 port map( A1 => n9652, A2 => n30274, B1 => n17816, B2 => 
                           n30268, ZN => n28901);
   U23197 : AOI221_X1 port map( B1 => n30286, B2 => n22200, C1 => n30280, C2 =>
                           n9715, A => n28882, ZN => n28877);
   U23198 : OAI22_X1 port map( A1 => n9651, A2 => n30274, B1 => n17815, B2 => 
                           n30268, ZN => n28882);
   U23199 : AOI221_X1 port map( B1 => n30286, B2 => n22201, C1 => n30280, C2 =>
                           n9714, A => n28863, ZN => n28858);
   U23200 : OAI22_X1 port map( A1 => n9650, A2 => n30274, B1 => n17814, B2 => 
                           n30268, ZN => n28863);
   U23201 : AOI221_X1 port map( B1 => n30286, B2 => n22202, C1 => n30280, C2 =>
                           n9713, A => n28844, ZN => n28839);
   U23202 : OAI22_X1 port map( A1 => n9649, A2 => n30274, B1 => n17813, B2 => 
                           n30268, ZN => n28844);
   U23203 : AOI221_X1 port map( B1 => n30287, B2 => n22203, C1 => n30281, C2 =>
                           n9712, A => n28825, ZN => n28820);
   U23204 : OAI22_X1 port map( A1 => n9648, A2 => n30275, B1 => n17812, B2 => 
                           n30269, ZN => n28825);
   U23205 : AOI221_X1 port map( B1 => n30287, B2 => n22204, C1 => n30281, C2 =>
                           n9711, A => n28806, ZN => n28801);
   U23206 : OAI22_X1 port map( A1 => n9647, A2 => n30275, B1 => n17811, B2 => 
                           n30269, ZN => n28806);
   U23207 : AOI221_X1 port map( B1 => n30287, B2 => n22205, C1 => n30281, C2 =>
                           n9710, A => n28787, ZN => n28782);
   U23208 : OAI22_X1 port map( A1 => n9646, A2 => n30275, B1 => n17810, B2 => 
                           n30269, ZN => n28787);
   U23209 : AOI221_X1 port map( B1 => n30287, B2 => n22206, C1 => n30281, C2 =>
                           n9709, A => n28768, ZN => n28763);
   U23210 : OAI22_X1 port map( A1 => n9645, A2 => n30275, B1 => n17809, B2 => 
                           n30269, ZN => n28768);
   U23211 : AOI221_X1 port map( B1 => n30287, B2 => n22207, C1 => n30281, C2 =>
                           n9708, A => n28749, ZN => n28744);
   U23212 : OAI22_X1 port map( A1 => n9644, A2 => n30275, B1 => n17808, B2 => 
                           n30269, ZN => n28749);
   U23213 : AOI221_X1 port map( B1 => n30287, B2 => n22208, C1 => n30281, C2 =>
                           n9707, A => n28730, ZN => n28725);
   U23214 : OAI22_X1 port map( A1 => n9643, A2 => n30275, B1 => n17807, B2 => 
                           n30269, ZN => n28730);
   U23215 : AOI221_X1 port map( B1 => n30287, B2 => n22209, C1 => n30281, C2 =>
                           n9706, A => n28711, ZN => n28706);
   U23216 : OAI22_X1 port map( A1 => n9642, A2 => n30275, B1 => n17806, B2 => 
                           n30269, ZN => n28711);
   U23217 : AOI221_X1 port map( B1 => n30287, B2 => n22210, C1 => n30281, C2 =>
                           n9705, A => n28692, ZN => n28687);
   U23218 : OAI22_X1 port map( A1 => n9641, A2 => n30275, B1 => n17805, B2 => 
                           n30269, ZN => n28692);
   U23219 : AOI221_X1 port map( B1 => n30287, B2 => n22211, C1 => n30281, C2 =>
                           n9704, A => n28673, ZN => n28668);
   U23220 : OAI22_X1 port map( A1 => n9640, A2 => n30275, B1 => n17804, B2 => 
                           n30269, ZN => n28673);
   U23221 : AOI221_X1 port map( B1 => n30287, B2 => n22212, C1 => n30281, C2 =>
                           n9703, A => n28654, ZN => n28649);
   U23222 : OAI22_X1 port map( A1 => n9639, A2 => n30275, B1 => n17803, B2 => 
                           n30269, ZN => n28654);
   U23223 : AOI221_X1 port map( B1 => n30287, B2 => n22213, C1 => n30281, C2 =>
                           n9702, A => n28635, ZN => n28630);
   U23224 : OAI22_X1 port map( A1 => n9638, A2 => n30275, B1 => n17802, B2 => 
                           n30269, ZN => n28635);
   U23225 : AOI221_X1 port map( B1 => n30287, B2 => n22214, C1 => n30281, C2 =>
                           n9701, A => n28616, ZN => n28611);
   U23226 : OAI22_X1 port map( A1 => n9637, A2 => n30275, B1 => n17801, B2 => 
                           n30269, ZN => n28616);
   U23227 : AOI221_X1 port map( B1 => n30288, B2 => n22215, C1 => n30282, C2 =>
                           n9700, A => n28597, ZN => n28592);
   U23228 : OAI22_X1 port map( A1 => n9636, A2 => n30276, B1 => n17800, B2 => 
                           n30270, ZN => n28597);
   U23229 : AOI221_X1 port map( B1 => n30288, B2 => n22216, C1 => n30282, C2 =>
                           n9699, A => n28578, ZN => n28573);
   U23230 : OAI22_X1 port map( A1 => n9635, A2 => n30276, B1 => n17799, B2 => 
                           n30270, ZN => n28578);
   U23231 : AOI221_X1 port map( B1 => n30288, B2 => n22217, C1 => n30282, C2 =>
                           n9698, A => n28559, ZN => n28554);
   U23232 : OAI22_X1 port map( A1 => n9634, A2 => n30276, B1 => n17798, B2 => 
                           n30270, ZN => n28559);
   U23233 : AOI221_X1 port map( B1 => n30288, B2 => n22218, C1 => n30282, C2 =>
                           n9697, A => n28540, ZN => n28535);
   U23234 : OAI22_X1 port map( A1 => n9633, A2 => n30276, B1 => n17797, B2 => 
                           n30270, ZN => n28540);
   U23235 : AOI221_X1 port map( B1 => n30288, B2 => n22219, C1 => n30282, C2 =>
                           n9696, A => n28521, ZN => n28516);
   U23236 : OAI22_X1 port map( A1 => n9632, A2 => n30276, B1 => n17796, B2 => 
                           n30270, ZN => n28521);
   U23237 : AOI221_X1 port map( B1 => n30288, B2 => n22220, C1 => n30282, C2 =>
                           n9695, A => n28502, ZN => n28497);
   U23238 : OAI22_X1 port map( A1 => n9631, A2 => n30276, B1 => n17795, B2 => 
                           n30270, ZN => n28502);
   U23239 : AOI221_X1 port map( B1 => n30288, B2 => n22221, C1 => n30282, C2 =>
                           n9694, A => n28483, ZN => n28478);
   U23240 : OAI22_X1 port map( A1 => n9630, A2 => n30276, B1 => n17794, B2 => 
                           n30270, ZN => n28483);
   U23241 : AOI221_X1 port map( B1 => n30288, B2 => n22222, C1 => n30282, C2 =>
                           n9693, A => n28464, ZN => n28459);
   U23242 : OAI22_X1 port map( A1 => n9629, A2 => n30276, B1 => n17793, B2 => 
                           n30270, ZN => n28464);
   U23243 : AOI221_X1 port map( B1 => n30288, B2 => n22223, C1 => n30282, C2 =>
                           n9692, A => n28445, ZN => n28440);
   U23244 : OAI22_X1 port map( A1 => n9628, A2 => n30276, B1 => n17792, B2 => 
                           n30270, ZN => n28445);
   U23245 : AOI221_X1 port map( B1 => n30288, B2 => n22224, C1 => n30282, C2 =>
                           n9691, A => n28426, ZN => n28421);
   U23246 : OAI22_X1 port map( A1 => n9627, A2 => n30276, B1 => n17791, B2 => 
                           n30270, ZN => n28426);
   U23247 : AOI221_X1 port map( B1 => n30288, B2 => n22225, C1 => n30282, C2 =>
                           n9690, A => n28407, ZN => n28402);
   U23248 : OAI22_X1 port map( A1 => n9626, A2 => n30276, B1 => n17790, B2 => 
                           n30270, ZN => n28407);
   U23249 : AOI221_X1 port map( B1 => n30288, B2 => n22226, C1 => n30282, C2 =>
                           n9689, A => n28388, ZN => n28383);
   U23250 : OAI22_X1 port map( A1 => n9625, A2 => n30276, B1 => n17789, B2 => 
                           n30270, ZN => n28388);
   U23251 : AOI221_X1 port map( B1 => n30289, B2 => n22227, C1 => n30283, C2 =>
                           n9688, A => n28369, ZN => n28364);
   U23252 : OAI22_X1 port map( A1 => n9624, A2 => n30277, B1 => n17788, B2 => 
                           n30271, ZN => n28369);
   U23253 : AOI221_X1 port map( B1 => n30289, B2 => n22228, C1 => n30283, C2 =>
                           n9687, A => n28350, ZN => n28345);
   U23254 : OAI22_X1 port map( A1 => n9623, A2 => n30277, B1 => n17787, B2 => 
                           n30271, ZN => n28350);
   U23255 : AOI221_X1 port map( B1 => n30289, B2 => n22229, C1 => n30283, C2 =>
                           n9686, A => n28331, ZN => n28326);
   U23256 : OAI22_X1 port map( A1 => n9622, A2 => n30277, B1 => n17786, B2 => 
                           n30271, ZN => n28331);
   U23257 : AOI221_X1 port map( B1 => n30289, B2 => n22230, C1 => n30283, C2 =>
                           n9685, A => n28312, ZN => n28307);
   U23258 : OAI22_X1 port map( A1 => n9621, A2 => n30277, B1 => n17785, B2 => 
                           n30271, ZN => n28312);
   U23259 : AOI221_X1 port map( B1 => n30289, B2 => n22231, C1 => n30283, C2 =>
                           n9684, A => n28293, ZN => n28288);
   U23260 : OAI22_X1 port map( A1 => n9620, A2 => n30277, B1 => n17784, B2 => 
                           n30271, ZN => n28293);
   U23261 : AOI221_X1 port map( B1 => n30289, B2 => n22232, C1 => n30283, C2 =>
                           n9683, A => n28274, ZN => n28269);
   U23262 : OAI22_X1 port map( A1 => n9619, A2 => n30277, B1 => n17783, B2 => 
                           n30271, ZN => n28274);
   U23263 : AOI221_X1 port map( B1 => n30289, B2 => n22233, C1 => n30283, C2 =>
                           n9682, A => n28255, ZN => n28250);
   U23264 : OAI22_X1 port map( A1 => n9618, A2 => n30277, B1 => n17782, B2 => 
                           n30271, ZN => n28255);
   U23265 : AOI221_X1 port map( B1 => n30289, B2 => n22234, C1 => n30283, C2 =>
                           n9681, A => n28236, ZN => n28231);
   U23266 : OAI22_X1 port map( A1 => n9617, A2 => n30277, B1 => n17781, B2 => 
                           n30271, ZN => n28236);
   U23267 : AOI221_X1 port map( B1 => n30289, B2 => n22235, C1 => n30283, C2 =>
                           n9680, A => n28217, ZN => n28212);
   U23268 : OAI22_X1 port map( A1 => n9616, A2 => n30277, B1 => n17780, B2 => 
                           n30271, ZN => n28217);
   U23269 : AOI221_X1 port map( B1 => n30289, B2 => n22236, C1 => n30283, C2 =>
                           n9679, A => n28198, ZN => n28193);
   U23270 : OAI22_X1 port map( A1 => n9615, A2 => n30277, B1 => n17779, B2 => 
                           n30271, ZN => n28198);
   U23271 : AOI221_X1 port map( B1 => n30289, B2 => n22237, C1 => n30283, C2 =>
                           n9678, A => n28179, ZN => n28174);
   U23272 : OAI22_X1 port map( A1 => n9614, A2 => n30277, B1 => n17778, B2 => 
                           n30271, ZN => n28179);
   U23273 : AOI221_X1 port map( B1 => n30289, B2 => n22238, C1 => n30283, C2 =>
                           n9677, A => n28160, ZN => n28155);
   U23274 : OAI22_X1 port map( A1 => n9613, A2 => n30277, B1 => n17777, B2 => 
                           n30271, ZN => n28160);
   U23275 : AOI221_X1 port map( B1 => n30333, B2 => n21806, C1 => n30327, C2 =>
                           n9549, A => n29070, ZN => n29069);
   U23276 : OAI22_X1 port map( A1 => n9229, A2 => n30321, B1 => n9997, B2 => 
                           n30315, ZN => n29070);
   U23277 : AOI221_X1 port map( B1 => n30334, B2 => n21807, C1 => n30328, C2 =>
                           n9544, A => n29051, ZN => n29050);
   U23278 : OAI22_X1 port map( A1 => n9224, A2 => n30322, B1 => n9992, B2 => 
                           n30316, ZN => n29051);
   U23279 : AOI221_X1 port map( B1 => n30334, B2 => n21808, C1 => n30328, C2 =>
                           n9539, A => n29032, ZN => n29031);
   U23280 : OAI22_X1 port map( A1 => n9219, A2 => n30322, B1 => n9987, B2 => 
                           n30316, ZN => n29032);
   U23281 : AOI221_X1 port map( B1 => n30334, B2 => n21809, C1 => n30328, C2 =>
                           n9534, A => n29013, ZN => n29012);
   U23282 : OAI22_X1 port map( A1 => n9214, A2 => n30322, B1 => n9982, B2 => 
                           n30316, ZN => n29013);
   U23283 : AOI221_X1 port map( B1 => n30334, B2 => n21810, C1 => n30328, C2 =>
                           n9529, A => n28994, ZN => n28993);
   U23284 : OAI22_X1 port map( A1 => n9209, A2 => n30322, B1 => n9977, B2 => 
                           n30316, ZN => n28994);
   U23285 : AOI221_X1 port map( B1 => n30334, B2 => n21811, C1 => n30328, C2 =>
                           n9524, A => n28975, ZN => n28974);
   U23286 : OAI22_X1 port map( A1 => n9204, A2 => n30322, B1 => n9972, B2 => 
                           n30316, ZN => n28975);
   U23287 : AOI221_X1 port map( B1 => n30334, B2 => n21812, C1 => n30328, C2 =>
                           n9519, A => n28956, ZN => n28955);
   U23288 : OAI22_X1 port map( A1 => n9199, A2 => n30322, B1 => n9967, B2 => 
                           n30316, ZN => n28956);
   U23289 : AOI221_X1 port map( B1 => n30334, B2 => n21813, C1 => n30328, C2 =>
                           n9514, A => n28937, ZN => n28936);
   U23290 : OAI22_X1 port map( A1 => n9194, A2 => n30322, B1 => n9962, B2 => 
                           n30316, ZN => n28937);
   U23291 : AOI221_X1 port map( B1 => n30334, B2 => n21814, C1 => n30328, C2 =>
                           n9509, A => n28918, ZN => n28917);
   U23292 : OAI22_X1 port map( A1 => n9189, A2 => n30322, B1 => n9957, B2 => 
                           n30316, ZN => n28918);
   U23293 : AOI221_X1 port map( B1 => n30334, B2 => n21815, C1 => n30328, C2 =>
                           n9504, A => n28899, ZN => n28898);
   U23294 : OAI22_X1 port map( A1 => n9184, A2 => n30322, B1 => n9952, B2 => 
                           n30316, ZN => n28899);
   U23295 : AOI221_X1 port map( B1 => n30334, B2 => n21816, C1 => n30328, C2 =>
                           n9499, A => n28880, ZN => n28879);
   U23296 : OAI22_X1 port map( A1 => n9179, A2 => n30322, B1 => n9947, B2 => 
                           n30316, ZN => n28880);
   U23297 : AOI221_X1 port map( B1 => n30334, B2 => n21817, C1 => n30328, C2 =>
                           n9494, A => n28861, ZN => n28860);
   U23298 : OAI22_X1 port map( A1 => n9174, A2 => n30322, B1 => n9942, B2 => 
                           n30316, ZN => n28861);
   U23299 : AOI221_X1 port map( B1 => n30334, B2 => n21818, C1 => n30328, C2 =>
                           n9489, A => n28842, ZN => n28841);
   U23300 : OAI22_X1 port map( A1 => n9169, A2 => n30322, B1 => n9937, B2 => 
                           n30316, ZN => n28842);
   U23301 : AOI221_X1 port map( B1 => n30335, B2 => n21819, C1 => n30329, C2 =>
                           n9484, A => n28823, ZN => n28822);
   U23302 : OAI22_X1 port map( A1 => n9164, A2 => n30323, B1 => n9932, B2 => 
                           n30317, ZN => n28823);
   U23303 : AOI221_X1 port map( B1 => n30335, B2 => n21820, C1 => n30329, C2 =>
                           n9479, A => n28804, ZN => n28803);
   U23304 : OAI22_X1 port map( A1 => n9159, A2 => n30323, B1 => n9927, B2 => 
                           n30317, ZN => n28804);
   U23305 : AOI221_X1 port map( B1 => n30335, B2 => n21821, C1 => n30329, C2 =>
                           n9474, A => n28785, ZN => n28784);
   U23306 : OAI22_X1 port map( A1 => n9154, A2 => n30323, B1 => n9922, B2 => 
                           n30317, ZN => n28785);
   U23307 : AOI221_X1 port map( B1 => n30335, B2 => n21822, C1 => n30329, C2 =>
                           n9469, A => n28766, ZN => n28765);
   U23308 : OAI22_X1 port map( A1 => n9149, A2 => n30323, B1 => n9917, B2 => 
                           n30317, ZN => n28766);
   U23309 : AOI221_X1 port map( B1 => n30335, B2 => n21823, C1 => n30329, C2 =>
                           n9464, A => n28747, ZN => n28746);
   U23310 : OAI22_X1 port map( A1 => n9144, A2 => n30323, B1 => n9912, B2 => 
                           n30317, ZN => n28747);
   U23311 : AOI221_X1 port map( B1 => n30335, B2 => n21824, C1 => n30329, C2 =>
                           n9459, A => n28728, ZN => n28727);
   U23312 : OAI22_X1 port map( A1 => n9139, A2 => n30323, B1 => n9907, B2 => 
                           n30317, ZN => n28728);
   U23313 : AOI221_X1 port map( B1 => n30335, B2 => n21825, C1 => n30329, C2 =>
                           n9454, A => n28709, ZN => n28708);
   U23314 : OAI22_X1 port map( A1 => n9134, A2 => n30323, B1 => n9902, B2 => 
                           n30317, ZN => n28709);
   U23315 : AOI221_X1 port map( B1 => n30335, B2 => n21826, C1 => n30329, C2 =>
                           n9449, A => n28690, ZN => n28689);
   U23316 : OAI22_X1 port map( A1 => n9129, A2 => n30323, B1 => n9897, B2 => 
                           n30317, ZN => n28690);
   U23317 : AOI221_X1 port map( B1 => n30335, B2 => n21827, C1 => n30329, C2 =>
                           n9444, A => n28671, ZN => n28670);
   U23318 : OAI22_X1 port map( A1 => n9124, A2 => n30323, B1 => n9892, B2 => 
                           n30317, ZN => n28671);
   U23319 : AOI221_X1 port map( B1 => n30335, B2 => n21828, C1 => n30329, C2 =>
                           n9439, A => n28652, ZN => n28651);
   U23320 : OAI22_X1 port map( A1 => n9119, A2 => n30323, B1 => n9887, B2 => 
                           n30317, ZN => n28652);
   U23321 : AOI221_X1 port map( B1 => n30335, B2 => n21829, C1 => n30329, C2 =>
                           n9434, A => n28633, ZN => n28632);
   U23322 : OAI22_X1 port map( A1 => n9114, A2 => n30323, B1 => n9882, B2 => 
                           n30317, ZN => n28633);
   U23323 : AOI221_X1 port map( B1 => n30335, B2 => n21830, C1 => n30329, C2 =>
                           n9429, A => n28614, ZN => n28613);
   U23324 : OAI22_X1 port map( A1 => n9109, A2 => n30323, B1 => n9877, B2 => 
                           n30317, ZN => n28614);
   U23325 : AOI221_X1 port map( B1 => n30336, B2 => n21831, C1 => n30330, C2 =>
                           n9424, A => n28595, ZN => n28594);
   U23326 : OAI22_X1 port map( A1 => n9104, A2 => n30324, B1 => n9872, B2 => 
                           n30318, ZN => n28595);
   U23327 : AOI221_X1 port map( B1 => n30336, B2 => n21832, C1 => n30330, C2 =>
                           n9419, A => n28576, ZN => n28575);
   U23328 : OAI22_X1 port map( A1 => n9099, A2 => n30324, B1 => n9867, B2 => 
                           n30318, ZN => n28576);
   U23329 : AOI221_X1 port map( B1 => n30336, B2 => n21833, C1 => n30330, C2 =>
                           n9414, A => n28557, ZN => n28556);
   U23330 : OAI22_X1 port map( A1 => n9094, A2 => n30324, B1 => n9862, B2 => 
                           n30318, ZN => n28557);
   U23331 : AOI221_X1 port map( B1 => n30336, B2 => n21834, C1 => n30330, C2 =>
                           n9409, A => n28538, ZN => n28537);
   U23332 : OAI22_X1 port map( A1 => n9089, A2 => n30324, B1 => n9857, B2 => 
                           n30318, ZN => n28538);
   U23333 : AOI221_X1 port map( B1 => n30336, B2 => n21835, C1 => n30330, C2 =>
                           n9404, A => n28519, ZN => n28518);
   U23334 : OAI22_X1 port map( A1 => n9084, A2 => n30324, B1 => n9852, B2 => 
                           n30318, ZN => n28519);
   U23335 : AOI221_X1 port map( B1 => n30336, B2 => n21836, C1 => n30330, C2 =>
                           n9399, A => n28500, ZN => n28499);
   U23336 : OAI22_X1 port map( A1 => n9079, A2 => n30324, B1 => n9847, B2 => 
                           n30318, ZN => n28500);
   U23337 : AOI221_X1 port map( B1 => n30336, B2 => n21837, C1 => n30330, C2 =>
                           n9394, A => n28481, ZN => n28480);
   U23338 : OAI22_X1 port map( A1 => n9074, A2 => n30324, B1 => n9842, B2 => 
                           n30318, ZN => n28481);
   U23339 : AOI221_X1 port map( B1 => n30336, B2 => n21838, C1 => n30330, C2 =>
                           n9389, A => n28462, ZN => n28461);
   U23340 : OAI22_X1 port map( A1 => n9069, A2 => n30324, B1 => n9837, B2 => 
                           n30318, ZN => n28462);
   U23341 : AOI221_X1 port map( B1 => n30336, B2 => n21839, C1 => n30330, C2 =>
                           n9384, A => n28443, ZN => n28442);
   U23342 : OAI22_X1 port map( A1 => n9064, A2 => n30324, B1 => n9832, B2 => 
                           n30318, ZN => n28443);
   U23343 : AOI221_X1 port map( B1 => n30336, B2 => n21840, C1 => n30330, C2 =>
                           n9379, A => n28424, ZN => n28423);
   U23344 : OAI22_X1 port map( A1 => n9059, A2 => n30324, B1 => n9827, B2 => 
                           n30318, ZN => n28424);
   U23345 : AOI221_X1 port map( B1 => n30336, B2 => n21841, C1 => n30330, C2 =>
                           n9374, A => n28405, ZN => n28404);
   U23346 : OAI22_X1 port map( A1 => n9054, A2 => n30324, B1 => n9822, B2 => 
                           n30318, ZN => n28405);
   U23347 : AOI221_X1 port map( B1 => n30336, B2 => n21842, C1 => n30330, C2 =>
                           n9369, A => n28386, ZN => n28385);
   U23348 : OAI22_X1 port map( A1 => n9049, A2 => n30324, B1 => n9817, B2 => 
                           n30318, ZN => n28386);
   U23349 : AOI221_X1 port map( B1 => n30337, B2 => n21843, C1 => n30331, C2 =>
                           n9364, A => n28367, ZN => n28366);
   U23350 : OAI22_X1 port map( A1 => n9044, A2 => n30325, B1 => n9812, B2 => 
                           n30319, ZN => n28367);
   U23351 : AOI221_X1 port map( B1 => n30337, B2 => n21844, C1 => n30331, C2 =>
                           n9359, A => n28348, ZN => n28347);
   U23352 : OAI22_X1 port map( A1 => n9039, A2 => n30325, B1 => n9807, B2 => 
                           n30319, ZN => n28348);
   U23353 : AOI221_X1 port map( B1 => n30337, B2 => n21845, C1 => n30331, C2 =>
                           n9354, A => n28329, ZN => n28328);
   U23354 : OAI22_X1 port map( A1 => n9034, A2 => n30325, B1 => n9802, B2 => 
                           n30319, ZN => n28329);
   U23355 : AOI221_X1 port map( B1 => n30337, B2 => n21846, C1 => n30331, C2 =>
                           n9349, A => n28310, ZN => n28309);
   U23356 : OAI22_X1 port map( A1 => n9029, A2 => n30325, B1 => n9797, B2 => 
                           n30319, ZN => n28310);
   U23357 : AOI221_X1 port map( B1 => n30337, B2 => n21847, C1 => n30331, C2 =>
                           n9344, A => n28291, ZN => n28290);
   U23358 : OAI22_X1 port map( A1 => n9024, A2 => n30325, B1 => n9792, B2 => 
                           n30319, ZN => n28291);
   U23359 : AOI221_X1 port map( B1 => n30337, B2 => n21848, C1 => n30331, C2 =>
                           n9339, A => n28272, ZN => n28271);
   U23360 : OAI22_X1 port map( A1 => n9019, A2 => n30325, B1 => n9787, B2 => 
                           n30319, ZN => n28272);
   U23361 : AOI221_X1 port map( B1 => n30337, B2 => n21849, C1 => n30331, C2 =>
                           n9334, A => n28253, ZN => n28252);
   U23362 : OAI22_X1 port map( A1 => n9014, A2 => n30325, B1 => n9782, B2 => 
                           n30319, ZN => n28253);
   U23363 : AOI221_X1 port map( B1 => n30337, B2 => n21850, C1 => n30331, C2 =>
                           n9329, A => n28234, ZN => n28233);
   U23364 : OAI22_X1 port map( A1 => n9009, A2 => n30325, B1 => n9777, B2 => 
                           n30319, ZN => n28234);
   U23365 : AOI221_X1 port map( B1 => n30337, B2 => n21851, C1 => n30331, C2 =>
                           n9324, A => n28215, ZN => n28214);
   U23366 : OAI22_X1 port map( A1 => n9004, A2 => n30325, B1 => n9772, B2 => 
                           n30319, ZN => n28215);
   U23367 : AOI221_X1 port map( B1 => n30337, B2 => n21852, C1 => n30331, C2 =>
                           n9319, A => n28196, ZN => n28195);
   U23368 : OAI22_X1 port map( A1 => n8999, A2 => n30325, B1 => n9767, B2 => 
                           n30319, ZN => n28196);
   U23369 : AOI221_X1 port map( B1 => n30337, B2 => n21853, C1 => n30331, C2 =>
                           n9314, A => n28177, ZN => n28176);
   U23370 : OAI22_X1 port map( A1 => n8994, A2 => n30325, B1 => n9762, B2 => 
                           n30319, ZN => n28177);
   U23371 : AOI221_X1 port map( B1 => n30337, B2 => n21854, C1 => n30331, C2 =>
                           n9309, A => n28158, ZN => n28157);
   U23372 : OAI22_X1 port map( A1 => n8989, A2 => n30325, B1 => n9757, B2 => 
                           n30319, ZN => n28158);
   U23373 : AOI221_X1 port map( B1 => n30213, B2 => n21859, C1 => n30207, C2 =>
                           n9608, A => n29301, ZN => n29296);
   U23374 : OAI22_X1 port map( A1 => n26088, A2 => n30201, B1 => n26022, B2 => 
                           n30195, ZN => n29301);
   U23375 : AOI221_X1 port map( B1 => n30333, B2 => n21795, C1 => n30327, C2 =>
                           n9604, A => n29280, ZN => n29279);
   U23376 : OAI22_X1 port map( A1 => n9284, A2 => n30321, B1 => n25229, B2 => 
                           n30315, ZN => n29280);
   U23377 : AOI221_X1 port map( B1 => n30213, B2 => n21860, C1 => n30207, C2 =>
                           n9603, A => n29269, ZN => n29266);
   U23378 : OAI22_X1 port map( A1 => n26087, A2 => n30201, B1 => n26021, B2 => 
                           n30195, ZN => n29269);
   U23379 : AOI221_X1 port map( B1 => n30333, B2 => n21796, C1 => n30327, C2 =>
                           n9599, A => n29260, ZN => n29259);
   U23380 : OAI22_X1 port map( A1 => n9279, A2 => n30321, B1 => n25227, B2 => 
                           n30315, ZN => n29260);
   U23381 : AOI221_X1 port map( B1 => n30213, B2 => n21861, C1 => n30207, C2 =>
                           n9598, A => n29250, ZN => n29247);
   U23382 : OAI22_X1 port map( A1 => n26086, A2 => n30201, B1 => n26020, B2 => 
                           n30195, ZN => n29250);
   U23383 : AOI221_X1 port map( B1 => n30333, B2 => n21797, C1 => n30327, C2 =>
                           n9594, A => n29241, ZN => n29240);
   U23384 : OAI22_X1 port map( A1 => n9274, A2 => n30321, B1 => n25225, B2 => 
                           n30315, ZN => n29241);
   U23385 : AOI221_X1 port map( B1 => n30213, B2 => n21862, C1 => n30207, C2 =>
                           n9593, A => n29231, ZN => n29228);
   U23386 : OAI22_X1 port map( A1 => n26085, A2 => n30201, B1 => n26019, B2 => 
                           n30195, ZN => n29231);
   U23387 : AOI221_X1 port map( B1 => n30333, B2 => n21798, C1 => n30327, C2 =>
                           n9589, A => n29222, ZN => n29221);
   U23388 : OAI22_X1 port map( A1 => n9269, A2 => n30321, B1 => n25223, B2 => 
                           n30315, ZN => n29222);
   U23389 : AOI221_X1 port map( B1 => n30213, B2 => n21863, C1 => n30207, C2 =>
                           n9588, A => n29212, ZN => n29209);
   U23390 : OAI22_X1 port map( A1 => n26084, A2 => n30201, B1 => n26018, B2 => 
                           n30195, ZN => n29212);
   U23391 : AOI221_X1 port map( B1 => n30333, B2 => n21799, C1 => n30327, C2 =>
                           n9584, A => n29203, ZN => n29202);
   U23392 : OAI22_X1 port map( A1 => n9264, A2 => n30321, B1 => n25221, B2 => 
                           n30315, ZN => n29203);
   U23393 : AOI221_X1 port map( B1 => n30213, B2 => n21864, C1 => n30207, C2 =>
                           n9583, A => n29193, ZN => n29190);
   U23394 : OAI22_X1 port map( A1 => n26083, A2 => n30201, B1 => n26017, B2 => 
                           n30195, ZN => n29193);
   U23395 : AOI221_X1 port map( B1 => n30333, B2 => n21800, C1 => n30327, C2 =>
                           n9579, A => n29184, ZN => n29183);
   U23396 : OAI22_X1 port map( A1 => n9259, A2 => n30321, B1 => n25219, B2 => 
                           n30315, ZN => n29184);
   U23397 : AOI221_X1 port map( B1 => n30213, B2 => n21865, C1 => n30207, C2 =>
                           n9578, A => n29174, ZN => n29171);
   U23398 : OAI22_X1 port map( A1 => n26082, A2 => n30201, B1 => n26016, B2 => 
                           n30195, ZN => n29174);
   U23399 : AOI221_X1 port map( B1 => n30333, B2 => n21801, C1 => n30327, C2 =>
                           n9574, A => n29165, ZN => n29164);
   U23400 : OAI22_X1 port map( A1 => n9254, A2 => n30321, B1 => n25217, B2 => 
                           n30315, ZN => n29165);
   U23401 : AOI221_X1 port map( B1 => n30213, B2 => n21866, C1 => n30207, C2 =>
                           n9573, A => n29155, ZN => n29152);
   U23402 : OAI22_X1 port map( A1 => n26081, A2 => n30201, B1 => n26015, B2 => 
                           n30195, ZN => n29155);
   U23403 : AOI221_X1 port map( B1 => n30333, B2 => n21802, C1 => n30327, C2 =>
                           n9569, A => n29146, ZN => n29145);
   U23404 : OAI22_X1 port map( A1 => n9249, A2 => n30321, B1 => n25215, B2 => 
                           n30315, ZN => n29146);
   U23405 : AOI221_X1 port map( B1 => n30213, B2 => n21867, C1 => n30207, C2 =>
                           n9568, A => n29136, ZN => n29133);
   U23406 : OAI22_X1 port map( A1 => n26080, A2 => n30201, B1 => n26014, B2 => 
                           n30195, ZN => n29136);
   U23407 : AOI221_X1 port map( B1 => n30333, B2 => n21803, C1 => n30327, C2 =>
                           n9564, A => n29127, ZN => n29126);
   U23408 : OAI22_X1 port map( A1 => n9244, A2 => n30321, B1 => n25213, B2 => 
                           n30315, ZN => n29127);
   U23409 : AOI221_X1 port map( B1 => n30213, B2 => n21868, C1 => n30207, C2 =>
                           n9563, A => n29117, ZN => n29114);
   U23410 : OAI22_X1 port map( A1 => n26079, A2 => n30201, B1 => n26013, B2 => 
                           n30195, ZN => n29117);
   U23411 : AOI221_X1 port map( B1 => n30333, B2 => n21804, C1 => n30327, C2 =>
                           n9559, A => n29108, ZN => n29107);
   U23412 : OAI22_X1 port map( A1 => n9239, A2 => n30321, B1 => n25211, B2 => 
                           n30315, ZN => n29108);
   U23413 : AOI221_X1 port map( B1 => n30213, B2 => n21869, C1 => n30207, C2 =>
                           n9558, A => n29098, ZN => n29095);
   U23414 : OAI22_X1 port map( A1 => n26078, A2 => n30201, B1 => n26012, B2 => 
                           n30195, ZN => n29098);
   U23415 : AOI221_X1 port map( B1 => n30333, B2 => n21805, C1 => n30327, C2 =>
                           n9554, A => n29089, ZN => n29088);
   U23416 : OAI22_X1 port map( A1 => n9234, A2 => n30321, B1 => n25209, B2 => 
                           n30315, ZN => n29089);
   U23417 : AOI221_X1 port map( B1 => n30213, B2 => n21870, C1 => n30207, C2 =>
                           n9553, A => n29079, ZN => n29076);
   U23418 : OAI22_X1 port map( A1 => n26077, A2 => n30201, B1 => n26011, B2 => 
                           n30195, ZN => n29079);
   U23419 : AOI221_X1 port map( B1 => n30214, B2 => n21871, C1 => n30208, C2 =>
                           n9548, A => n29060, ZN => n29057);
   U23420 : OAI22_X1 port map( A1 => n26076, A2 => n30202, B1 => n26010, B2 => 
                           n30196, ZN => n29060);
   U23421 : AOI221_X1 port map( B1 => n30214, B2 => n21872, C1 => n30208, C2 =>
                           n9543, A => n29041, ZN => n29038);
   U23422 : OAI22_X1 port map( A1 => n26075, A2 => n30202, B1 => n26009, B2 => 
                           n30196, ZN => n29041);
   U23423 : AOI221_X1 port map( B1 => n30214, B2 => n21873, C1 => n30208, C2 =>
                           n9538, A => n29022, ZN => n29019);
   U23424 : OAI22_X1 port map( A1 => n26074, A2 => n30202, B1 => n26008, B2 => 
                           n30196, ZN => n29022);
   U23425 : AOI221_X1 port map( B1 => n30214, B2 => n21874, C1 => n30208, C2 =>
                           n9533, A => n29003, ZN => n29000);
   U23426 : OAI22_X1 port map( A1 => n26073, A2 => n30202, B1 => n26007, B2 => 
                           n30196, ZN => n29003);
   U23427 : AOI221_X1 port map( B1 => n30214, B2 => n21875, C1 => n30208, C2 =>
                           n9528, A => n28984, ZN => n28981);
   U23428 : OAI22_X1 port map( A1 => n26072, A2 => n30202, B1 => n26006, B2 => 
                           n30196, ZN => n28984);
   U23429 : AOI221_X1 port map( B1 => n30214, B2 => n21876, C1 => n30208, C2 =>
                           n9523, A => n28965, ZN => n28962);
   U23430 : OAI22_X1 port map( A1 => n26071, A2 => n30202, B1 => n26005, B2 => 
                           n30196, ZN => n28965);
   U23431 : AOI221_X1 port map( B1 => n30214, B2 => n21877, C1 => n30208, C2 =>
                           n9518, A => n28946, ZN => n28943);
   U23432 : OAI22_X1 port map( A1 => n26070, A2 => n30202, B1 => n26004, B2 => 
                           n30196, ZN => n28946);
   U23433 : AOI221_X1 port map( B1 => n30214, B2 => n21878, C1 => n30208, C2 =>
                           n9513, A => n28927, ZN => n28924);
   U23434 : OAI22_X1 port map( A1 => n26069, A2 => n30202, B1 => n26003, B2 => 
                           n30196, ZN => n28927);
   U23435 : AOI221_X1 port map( B1 => n30214, B2 => n21879, C1 => n30208, C2 =>
                           n9508, A => n28908, ZN => n28905);
   U23436 : OAI22_X1 port map( A1 => n26068, A2 => n30202, B1 => n26002, B2 => 
                           n30196, ZN => n28908);
   U23437 : AOI221_X1 port map( B1 => n30214, B2 => n21880, C1 => n30208, C2 =>
                           n9503, A => n28889, ZN => n28886);
   U23438 : OAI22_X1 port map( A1 => n26067, A2 => n30202, B1 => n26001, B2 => 
                           n30196, ZN => n28889);
   U23439 : AOI221_X1 port map( B1 => n30214, B2 => n21881, C1 => n30208, C2 =>
                           n9498, A => n28870, ZN => n28867);
   U23440 : OAI22_X1 port map( A1 => n26066, A2 => n30202, B1 => n26000, B2 => 
                           n30196, ZN => n28870);
   U23441 : AOI221_X1 port map( B1 => n30214, B2 => n21882, C1 => n30208, C2 =>
                           n9493, A => n28851, ZN => n28848);
   U23442 : OAI22_X1 port map( A1 => n26065, A2 => n30202, B1 => n25999, B2 => 
                           n30196, ZN => n28851);
   U23443 : AOI221_X1 port map( B1 => n30215, B2 => n21883, C1 => n30209, C2 =>
                           n9488, A => n28832, ZN => n28829);
   U23444 : OAI22_X1 port map( A1 => n26064, A2 => n30203, B1 => n25998, B2 => 
                           n30197, ZN => n28832);
   U23445 : AOI221_X1 port map( B1 => n30215, B2 => n21884, C1 => n30209, C2 =>
                           n9483, A => n28813, ZN => n28810);
   U23446 : OAI22_X1 port map( A1 => n26063, A2 => n30203, B1 => n25997, B2 => 
                           n30197, ZN => n28813);
   U23447 : AOI221_X1 port map( B1 => n30215, B2 => n21885, C1 => n30209, C2 =>
                           n9478, A => n28794, ZN => n28791);
   U23448 : OAI22_X1 port map( A1 => n26062, A2 => n30203, B1 => n25996, B2 => 
                           n30197, ZN => n28794);
   U23449 : AOI221_X1 port map( B1 => n30215, B2 => n21886, C1 => n30209, C2 =>
                           n9473, A => n28775, ZN => n28772);
   U23450 : OAI22_X1 port map( A1 => n26061, A2 => n30203, B1 => n25995, B2 => 
                           n30197, ZN => n28775);
   U23451 : AOI221_X1 port map( B1 => n30215, B2 => n21887, C1 => n30209, C2 =>
                           n9468, A => n28756, ZN => n28753);
   U23452 : OAI22_X1 port map( A1 => n26060, A2 => n30203, B1 => n25994, B2 => 
                           n30197, ZN => n28756);
   U23453 : AOI221_X1 port map( B1 => n30215, B2 => n21888, C1 => n30209, C2 =>
                           n9463, A => n28737, ZN => n28734);
   U23454 : OAI22_X1 port map( A1 => n26059, A2 => n30203, B1 => n25993, B2 => 
                           n30197, ZN => n28737);
   U23455 : AOI221_X1 port map( B1 => n30215, B2 => n21889, C1 => n30209, C2 =>
                           n9458, A => n28718, ZN => n28715);
   U23456 : OAI22_X1 port map( A1 => n26058, A2 => n30203, B1 => n25992, B2 => 
                           n30197, ZN => n28718);
   U23457 : AOI221_X1 port map( B1 => n30215, B2 => n21890, C1 => n30209, C2 =>
                           n9453, A => n28699, ZN => n28696);
   U23458 : OAI22_X1 port map( A1 => n26057, A2 => n30203, B1 => n25991, B2 => 
                           n30197, ZN => n28699);
   U23459 : AOI221_X1 port map( B1 => n30215, B2 => n21891, C1 => n30209, C2 =>
                           n9448, A => n28680, ZN => n28677);
   U23460 : OAI22_X1 port map( A1 => n26056, A2 => n30203, B1 => n25990, B2 => 
                           n30197, ZN => n28680);
   U23461 : AOI221_X1 port map( B1 => n30215, B2 => n21892, C1 => n30209, C2 =>
                           n9443, A => n28661, ZN => n28658);
   U23462 : OAI22_X1 port map( A1 => n26055, A2 => n30203, B1 => n25989, B2 => 
                           n30197, ZN => n28661);
   U23463 : AOI221_X1 port map( B1 => n30215, B2 => n21893, C1 => n30209, C2 =>
                           n9438, A => n28642, ZN => n28639);
   U23464 : OAI22_X1 port map( A1 => n26054, A2 => n30203, B1 => n25988, B2 => 
                           n30197, ZN => n28642);
   U23465 : AOI221_X1 port map( B1 => n30215, B2 => n21894, C1 => n30209, C2 =>
                           n9433, A => n28623, ZN => n28620);
   U23466 : OAI22_X1 port map( A1 => n26053, A2 => n30203, B1 => n25987, B2 => 
                           n30197, ZN => n28623);
   U23467 : AOI221_X1 port map( B1 => n30216, B2 => n21895, C1 => n30210, C2 =>
                           n9428, A => n28604, ZN => n28601);
   U23468 : OAI22_X1 port map( A1 => n26052, A2 => n30204, B1 => n25986, B2 => 
                           n30198, ZN => n28604);
   U23469 : AOI221_X1 port map( B1 => n30216, B2 => n21896, C1 => n30210, C2 =>
                           n9423, A => n28585, ZN => n28582);
   U23470 : OAI22_X1 port map( A1 => n26051, A2 => n30204, B1 => n25985, B2 => 
                           n30198, ZN => n28585);
   U23471 : AOI221_X1 port map( B1 => n30216, B2 => n21897, C1 => n30210, C2 =>
                           n9418, A => n28566, ZN => n28563);
   U23472 : OAI22_X1 port map( A1 => n26050, A2 => n30204, B1 => n25984, B2 => 
                           n30198, ZN => n28566);
   U23473 : AOI221_X1 port map( B1 => n30216, B2 => n21898, C1 => n30210, C2 =>
                           n9413, A => n28547, ZN => n28544);
   U23474 : OAI22_X1 port map( A1 => n26049, A2 => n30204, B1 => n25983, B2 => 
                           n30198, ZN => n28547);
   U23475 : AOI221_X1 port map( B1 => n30216, B2 => n21899, C1 => n30210, C2 =>
                           n9408, A => n28528, ZN => n28525);
   U23476 : OAI22_X1 port map( A1 => n26048, A2 => n30204, B1 => n25982, B2 => 
                           n30198, ZN => n28528);
   U23477 : AOI221_X1 port map( B1 => n30216, B2 => n21900, C1 => n30210, C2 =>
                           n9403, A => n28509, ZN => n28506);
   U23478 : OAI22_X1 port map( A1 => n26047, A2 => n30204, B1 => n25981, B2 => 
                           n30198, ZN => n28509);
   U23479 : AOI221_X1 port map( B1 => n30216, B2 => n21901, C1 => n30210, C2 =>
                           n9398, A => n28490, ZN => n28487);
   U23480 : OAI22_X1 port map( A1 => n26046, A2 => n30204, B1 => n25980, B2 => 
                           n30198, ZN => n28490);
   U23481 : AOI221_X1 port map( B1 => n30216, B2 => n21902, C1 => n30210, C2 =>
                           n9393, A => n28471, ZN => n28468);
   U23482 : OAI22_X1 port map( A1 => n26045, A2 => n30204, B1 => n25979, B2 => 
                           n30198, ZN => n28471);
   U23483 : AOI221_X1 port map( B1 => n30216, B2 => n21903, C1 => n30210, C2 =>
                           n9388, A => n28452, ZN => n28449);
   U23484 : OAI22_X1 port map( A1 => n26044, A2 => n30204, B1 => n25978, B2 => 
                           n30198, ZN => n28452);
   U23485 : AOI221_X1 port map( B1 => n30216, B2 => n21904, C1 => n30210, C2 =>
                           n9383, A => n28433, ZN => n28430);
   U23486 : OAI22_X1 port map( A1 => n26043, A2 => n30204, B1 => n25977, B2 => 
                           n30198, ZN => n28433);
   U23487 : AOI221_X1 port map( B1 => n30216, B2 => n21905, C1 => n30210, C2 =>
                           n9378, A => n28414, ZN => n28411);
   U23488 : OAI22_X1 port map( A1 => n26042, A2 => n30204, B1 => n25976, B2 => 
                           n30198, ZN => n28414);
   U23489 : AOI221_X1 port map( B1 => n30216, B2 => n21906, C1 => n30210, C2 =>
                           n9373, A => n28395, ZN => n28392);
   U23490 : OAI22_X1 port map( A1 => n26041, A2 => n30204, B1 => n25975, B2 => 
                           n30198, ZN => n28395);
   U23491 : AOI221_X1 port map( B1 => n30217, B2 => n21907, C1 => n30211, C2 =>
                           n9368, A => n28376, ZN => n28373);
   U23492 : OAI22_X1 port map( A1 => n26040, A2 => n30205, B1 => n25974, B2 => 
                           n30199, ZN => n28376);
   U23493 : AOI221_X1 port map( B1 => n30217, B2 => n21908, C1 => n30211, C2 =>
                           n9363, A => n28357, ZN => n28354);
   U23494 : OAI22_X1 port map( A1 => n26039, A2 => n30205, B1 => n25973, B2 => 
                           n30199, ZN => n28357);
   U23495 : AOI221_X1 port map( B1 => n30217, B2 => n21909, C1 => n30211, C2 =>
                           n9358, A => n28338, ZN => n28335);
   U23496 : OAI22_X1 port map( A1 => n26038, A2 => n30205, B1 => n25972, B2 => 
                           n30199, ZN => n28338);
   U23497 : AOI221_X1 port map( B1 => n30217, B2 => n21910, C1 => n30211, C2 =>
                           n9353, A => n28319, ZN => n28316);
   U23498 : OAI22_X1 port map( A1 => n26037, A2 => n30205, B1 => n25971, B2 => 
                           n30199, ZN => n28319);
   U23499 : AOI221_X1 port map( B1 => n30217, B2 => n21911, C1 => n30211, C2 =>
                           n9348, A => n28300, ZN => n28297);
   U23500 : OAI22_X1 port map( A1 => n26036, A2 => n30205, B1 => n25970, B2 => 
                           n30199, ZN => n28300);
   U23501 : AOI221_X1 port map( B1 => n30217, B2 => n21912, C1 => n30211, C2 =>
                           n9343, A => n28281, ZN => n28278);
   U23502 : OAI22_X1 port map( A1 => n26035, A2 => n30205, B1 => n25969, B2 => 
                           n30199, ZN => n28281);
   U23503 : AOI221_X1 port map( B1 => n30217, B2 => n21913, C1 => n30211, C2 =>
                           n9338, A => n28262, ZN => n28259);
   U23504 : OAI22_X1 port map( A1 => n26034, A2 => n30205, B1 => n25968, B2 => 
                           n30199, ZN => n28262);
   U23505 : AOI221_X1 port map( B1 => n30217, B2 => n21914, C1 => n30211, C2 =>
                           n9333, A => n28243, ZN => n28240);
   U23506 : OAI22_X1 port map( A1 => n26033, A2 => n30205, B1 => n25967, B2 => 
                           n30199, ZN => n28243);
   U23507 : AOI221_X1 port map( B1 => n30217, B2 => n21915, C1 => n30211, C2 =>
                           n9328, A => n28224, ZN => n28221);
   U23508 : OAI22_X1 port map( A1 => n26032, A2 => n30205, B1 => n25966, B2 => 
                           n30199, ZN => n28224);
   U23509 : AOI221_X1 port map( B1 => n30217, B2 => n21916, C1 => n30211, C2 =>
                           n9323, A => n28205, ZN => n28202);
   U23510 : OAI22_X1 port map( A1 => n26031, A2 => n30205, B1 => n25965, B2 => 
                           n30199, ZN => n28205);
   U23511 : AOI221_X1 port map( B1 => n30217, B2 => n21917, C1 => n30211, C2 =>
                           n9318, A => n28186, ZN => n28183);
   U23512 : OAI22_X1 port map( A1 => n26030, A2 => n30205, B1 => n25964, B2 => 
                           n30199, ZN => n28186);
   U23513 : AOI221_X1 port map( B1 => n30217, B2 => n21918, C1 => n30211, C2 =>
                           n9313, A => n28167, ZN => n28164);
   U23514 : OAI22_X1 port map( A1 => n26029, A2 => n30205, B1 => n25963, B2 => 
                           n30199, ZN => n28167);
   U23515 : AOI221_X1 port map( B1 => n30468, B2 => n22089, C1 => n30462, C2 =>
                           n9482, A => n27351, ZN => n27344);
   U23516 : OAI22_X1 port map( A1 => n30457, A2 => n27340, B1 => n26290, B2 => 
                           n30449, ZN => n27351);
   U23517 : AOI221_X1 port map( B1 => n30468, B2 => n22090, C1 => n30462, C2 =>
                           n9477, A => n27325, ZN => n27318);
   U23518 : OAI22_X1 port map( A1 => n30457, A2 => n27314, B1 => n26289, B2 => 
                           n30449, ZN => n27325);
   U23519 : AOI221_X1 port map( B1 => n30468, B2 => n22091, C1 => n30462, C2 =>
                           n9472, A => n27299, ZN => n27292);
   U23520 : OAI22_X1 port map( A1 => n30457, A2 => n27288, B1 => n26288, B2 => 
                           n30449, ZN => n27299);
   U23521 : AOI221_X1 port map( B1 => n30468, B2 => n22092, C1 => n30462, C2 =>
                           n9467, A => n27273, ZN => n27266);
   U23522 : OAI22_X1 port map( A1 => n30457, A2 => n27262, B1 => n26287, B2 => 
                           n30449, ZN => n27273);
   U23523 : AOI221_X1 port map( B1 => n30468, B2 => n22093, C1 => n30462, C2 =>
                           n9462, A => n27247, ZN => n27240);
   U23524 : OAI22_X1 port map( A1 => n30457, A2 => n27236, B1 => n26286, B2 => 
                           n30449, ZN => n27247);
   U23525 : AOI221_X1 port map( B1 => n30468, B2 => n22094, C1 => n30462, C2 =>
                           n9457, A => n27221, ZN => n27214);
   U23526 : OAI22_X1 port map( A1 => n30457, A2 => n27210, B1 => n26285, B2 => 
                           n30449, ZN => n27221);
   U23527 : AOI221_X1 port map( B1 => n30468, B2 => n22095, C1 => n30462, C2 =>
                           n9452, A => n27195, ZN => n27188);
   U23528 : OAI22_X1 port map( A1 => n30457, A2 => n27184, B1 => n26284, B2 => 
                           n30449, ZN => n27195);
   U23529 : AOI221_X1 port map( B1 => n30468, B2 => n22096, C1 => n30462, C2 =>
                           n9447, A => n27169, ZN => n27162);
   U23530 : OAI22_X1 port map( A1 => n30457, A2 => n27158, B1 => n26283, B2 => 
                           n30449, ZN => n27169);
   U23531 : AOI221_X1 port map( B1 => n30468, B2 => n22097, C1 => n30462, C2 =>
                           n9442, A => n27143, ZN => n27136);
   U23532 : OAI22_X1 port map( A1 => n30457, A2 => n27132, B1 => n26282, B2 => 
                           n30449, ZN => n27143);
   U23533 : AOI221_X1 port map( B1 => n30468, B2 => n22098, C1 => n30462, C2 =>
                           n9437, A => n27117, ZN => n27110);
   U23534 : OAI22_X1 port map( A1 => n30457, A2 => n27106, B1 => n26281, B2 => 
                           n30449, ZN => n27117);
   U23535 : AOI221_X1 port map( B1 => n30468, B2 => n22099, C1 => n30462, C2 =>
                           n9432, A => n27091, ZN => n27084);
   U23536 : OAI22_X1 port map( A1 => n30457, A2 => n27080, B1 => n26280, B2 => 
                           n30449, ZN => n27091);
   U23537 : AOI221_X1 port map( B1 => n30469, B2 => n22100, C1 => n30463, C2 =>
                           n9427, A => n27065, ZN => n27058);
   U23538 : OAI22_X1 port map( A1 => n30457, A2 => n27054, B1 => n26279, B2 => 
                           n30450, ZN => n27065);
   U23539 : AOI221_X1 port map( B1 => n30469, B2 => n22101, C1 => n30463, C2 =>
                           n9422, A => n27039, ZN => n27032);
   U23540 : OAI22_X1 port map( A1 => n30457, A2 => n27028, B1 => n26278, B2 => 
                           n30450, ZN => n27039);
   U23541 : AOI221_X1 port map( B1 => n30469, B2 => n22102, C1 => n30463, C2 =>
                           n9417, A => n27013, ZN => n27006);
   U23542 : OAI22_X1 port map( A1 => n30456, A2 => n27002, B1 => n26277, B2 => 
                           n30450, ZN => n27013);
   U23543 : AOI221_X1 port map( B1 => n30469, B2 => n22103, C1 => n30463, C2 =>
                           n9412, A => n26987, ZN => n26980);
   U23544 : OAI22_X1 port map( A1 => n30456, A2 => n26976, B1 => n26276, B2 => 
                           n30450, ZN => n26987);
   U23545 : AOI221_X1 port map( B1 => n30469, B2 => n22104, C1 => n30463, C2 =>
                           n9407, A => n26961, ZN => n26954);
   U23546 : OAI22_X1 port map( A1 => n30456, A2 => n26950, B1 => n26275, B2 => 
                           n30450, ZN => n26961);
   U23547 : AOI221_X1 port map( B1 => n30469, B2 => n22105, C1 => n30463, C2 =>
                           n9402, A => n26935, ZN => n26928);
   U23548 : OAI22_X1 port map( A1 => n30456, A2 => n26924, B1 => n26274, B2 => 
                           n30450, ZN => n26935);
   U23549 : AOI221_X1 port map( B1 => n30469, B2 => n22106, C1 => n30463, C2 =>
                           n9397, A => n26909, ZN => n26902);
   U23550 : OAI22_X1 port map( A1 => n30456, A2 => n26898, B1 => n26273, B2 => 
                           n30450, ZN => n26909);
   U23551 : AOI221_X1 port map( B1 => n30469, B2 => n22107, C1 => n30463, C2 =>
                           n9392, A => n26883, ZN => n26876);
   U23552 : OAI22_X1 port map( A1 => n30456, A2 => n26872, B1 => n26272, B2 => 
                           n30450, ZN => n26883);
   U23553 : AOI221_X1 port map( B1 => n30469, B2 => n22108, C1 => n30463, C2 =>
                           n9387, A => n26857, ZN => n26850);
   U23554 : OAI22_X1 port map( A1 => n30456, A2 => n26846, B1 => n26271, B2 => 
                           n30450, ZN => n26857);
   U23555 : AOI221_X1 port map( B1 => n30469, B2 => n22109, C1 => n30463, C2 =>
                           n9382, A => n26831, ZN => n26824);
   U23556 : OAI22_X1 port map( A1 => n30456, A2 => n26820, B1 => n26270, B2 => 
                           n30450, ZN => n26831);
   U23557 : AOI221_X1 port map( B1 => n30469, B2 => n22110, C1 => n30463, C2 =>
                           n9377, A => n26805, ZN => n26798);
   U23558 : OAI22_X1 port map( A1 => n30456, A2 => n26794, B1 => n26269, B2 => 
                           n30450, ZN => n26805);
   U23559 : AOI221_X1 port map( B1 => n30469, B2 => n22111, C1 => n30463, C2 =>
                           n9372, A => n26779, ZN => n26772);
   U23560 : OAI22_X1 port map( A1 => n30456, A2 => n26768, B1 => n26268, B2 => 
                           n30450, ZN => n26779);
   U23561 : AOI221_X1 port map( B1 => n30470, B2 => n22112, C1 => n30464, C2 =>
                           n9367, A => n26753, ZN => n26746);
   U23562 : OAI22_X1 port map( A1 => n30456, A2 => n26742, B1 => n26267, B2 => 
                           n30451, ZN => n26753);
   U23563 : AOI221_X1 port map( B1 => n30470, B2 => n22113, C1 => n30464, C2 =>
                           n9362, A => n26727, ZN => n26720);
   U23564 : OAI22_X1 port map( A1 => n30456, A2 => n26716, B1 => n26266, B2 => 
                           n30451, ZN => n26727);
   U23565 : AOI221_X1 port map( B1 => n30470, B2 => n22114, C1 => n30464, C2 =>
                           n9357, A => n26701, ZN => n26694);
   U23566 : OAI22_X1 port map( A1 => n30456, A2 => n26690, B1 => n26265, B2 => 
                           n30451, ZN => n26701);
   U23567 : OAI22_X1 port map( A1 => n9992, A2 => n31146, B1 => n31137, B2 => 
                           n30980, ZN => n7829);
   U23568 : OAI22_X1 port map( A1 => n9987, A2 => n31146, B1 => n31137, B2 => 
                           n30983, ZN => n7830);
   U23569 : OAI22_X1 port map( A1 => n9982, A2 => n31146, B1 => n31137, B2 => 
                           n30986, ZN => n7831);
   U23570 : OAI22_X1 port map( A1 => n9977, A2 => n31146, B1 => n31137, B2 => 
                           n30989, ZN => n7832);
   U23571 : OAI22_X1 port map( A1 => n9972, A2 => n31146, B1 => n31137, B2 => 
                           n30992, ZN => n7833);
   U23572 : OAI22_X1 port map( A1 => n9967, A2 => n31145, B1 => n31137, B2 => 
                           n30995, ZN => n7834);
   U23573 : OAI22_X1 port map( A1 => n9962, A2 => n31145, B1 => n31137, B2 => 
                           n30998, ZN => n7835);
   U23574 : OAI22_X1 port map( A1 => n9957, A2 => n31145, B1 => n31137, B2 => 
                           n31001, ZN => n7836);
   U23575 : OAI22_X1 port map( A1 => n9952, A2 => n31145, B1 => n31137, B2 => 
                           n31004, ZN => n7837);
   U23576 : OAI22_X1 port map( A1 => n9947, A2 => n31145, B1 => n31137, B2 => 
                           n31007, ZN => n7838);
   U23577 : OAI22_X1 port map( A1 => n9942, A2 => n31145, B1 => n31137, B2 => 
                           n31010, ZN => n7839);
   U23578 : OAI22_X1 port map( A1 => n9937, A2 => n31145, B1 => n31137, B2 => 
                           n31013, ZN => n7840);
   U23579 : OAI22_X1 port map( A1 => n9932, A2 => n31145, B1 => n31138, B2 => 
                           n31016, ZN => n7841);
   U23580 : OAI22_X1 port map( A1 => n9927, A2 => n31145, B1 => n31138, B2 => 
                           n31019, ZN => n7842);
   U23581 : OAI22_X1 port map( A1 => n9922, A2 => n31145, B1 => n31138, B2 => 
                           n31022, ZN => n7843);
   U23582 : OAI22_X1 port map( A1 => n9917, A2 => n31145, B1 => n31138, B2 => 
                           n31025, ZN => n7844);
   U23583 : OAI22_X1 port map( A1 => n9912, A2 => n31145, B1 => n31138, B2 => 
                           n31028, ZN => n7845);
   U23584 : OAI22_X1 port map( A1 => n9907, A2 => n31144, B1 => n31138, B2 => 
                           n31031, ZN => n7846);
   U23585 : OAI22_X1 port map( A1 => n9902, A2 => n31144, B1 => n31138, B2 => 
                           n31034, ZN => n7847);
   U23586 : OAI22_X1 port map( A1 => n9897, A2 => n31144, B1 => n31138, B2 => 
                           n31037, ZN => n7848);
   U23587 : OAI22_X1 port map( A1 => n9892, A2 => n31144, B1 => n31138, B2 => 
                           n31040, ZN => n7849);
   U23588 : OAI22_X1 port map( A1 => n9887, A2 => n31144, B1 => n31138, B2 => 
                           n31043, ZN => n7850);
   U23589 : OAI22_X1 port map( A1 => n9882, A2 => n31144, B1 => n31138, B2 => 
                           n31046, ZN => n7851);
   U23590 : OAI22_X1 port map( A1 => n9877, A2 => n31144, B1 => n31138, B2 => 
                           n31049, ZN => n7852);
   U23591 : OAI22_X1 port map( A1 => n9872, A2 => n31144, B1 => n31139, B2 => 
                           n31052, ZN => n7853);
   U23592 : OAI22_X1 port map( A1 => n9867, A2 => n31144, B1 => n31139, B2 => 
                           n31055, ZN => n7854);
   U23593 : OAI22_X1 port map( A1 => n9862, A2 => n31144, B1 => n31139, B2 => 
                           n31058, ZN => n7855);
   U23594 : OAI22_X1 port map( A1 => n9857, A2 => n31144, B1 => n31139, B2 => 
                           n31061, ZN => n7856);
   U23595 : OAI22_X1 port map( A1 => n9852, A2 => n31143, B1 => n31139, B2 => 
                           n31064, ZN => n7857);
   U23596 : OAI22_X1 port map( A1 => n9847, A2 => n31143, B1 => n31139, B2 => 
                           n31067, ZN => n7858);
   U23597 : OAI22_X1 port map( A1 => n9842, A2 => n31143, B1 => n31139, B2 => 
                           n31070, ZN => n7859);
   U23598 : OAI22_X1 port map( A1 => n9837, A2 => n31143, B1 => n31139, B2 => 
                           n31073, ZN => n7860);
   U23599 : OAI22_X1 port map( A1 => n9832, A2 => n31143, B1 => n31139, B2 => 
                           n31076, ZN => n7861);
   U23600 : OAI22_X1 port map( A1 => n9827, A2 => n31143, B1 => n31139, B2 => 
                           n31079, ZN => n7862);
   U23601 : OAI22_X1 port map( A1 => n9822, A2 => n31143, B1 => n31139, B2 => 
                           n31082, ZN => n7863);
   U23602 : OAI22_X1 port map( A1 => n9817, A2 => n31143, B1 => n31139, B2 => 
                           n31085, ZN => n7864);
   U23603 : OAI22_X1 port map( A1 => n9812, A2 => n31143, B1 => n31140, B2 => 
                           n31088, ZN => n7865);
   U23604 : OAI22_X1 port map( A1 => n9807, A2 => n31143, B1 => n31140, B2 => 
                           n31091, ZN => n7866);
   U23605 : OAI22_X1 port map( A1 => n9802, A2 => n31143, B1 => n31140, B2 => 
                           n31094, ZN => n7867);
   U23606 : OAI22_X1 port map( A1 => n9797, A2 => n31143, B1 => n31140, B2 => 
                           n31097, ZN => n7868);
   U23607 : OAI22_X1 port map( A1 => n9792, A2 => n31142, B1 => n31140, B2 => 
                           n31100, ZN => n7869);
   U23608 : OAI22_X1 port map( A1 => n9787, A2 => n31142, B1 => n31140, B2 => 
                           n31103, ZN => n7870);
   U23609 : OAI22_X1 port map( A1 => n9782, A2 => n31142, B1 => n31140, B2 => 
                           n31106, ZN => n7871);
   U23610 : OAI22_X1 port map( A1 => n9777, A2 => n31142, B1 => n31140, B2 => 
                           n31109, ZN => n7872);
   U23611 : OAI22_X1 port map( A1 => n9772, A2 => n31142, B1 => n31140, B2 => 
                           n31112, ZN => n7873);
   U23612 : OAI22_X1 port map( A1 => n9767, A2 => n31142, B1 => n31140, B2 => 
                           n31115, ZN => n7874);
   U23613 : OAI22_X1 port map( A1 => n9762, A2 => n31142, B1 => n31140, B2 => 
                           n31118, ZN => n7875);
   U23614 : OAI22_X1 port map( A1 => n9757, A2 => n31142, B1 => n31140, B2 => 
                           n31121, ZN => n7876);
   U23615 : OAI22_X1 port map( A1 => n9752, A2 => n31142, B1 => n31141, B2 => 
                           n31124, ZN => n7877);
   U23616 : OAI22_X1 port map( A1 => n9747, A2 => n31142, B1 => n31141, B2 => 
                           n31127, ZN => n7878);
   U23617 : OAI22_X1 port map( A1 => n9742, A2 => n31142, B1 => n31141, B2 => 
                           n31130, ZN => n7879);
   U23618 : OAI22_X1 port map( A1 => n9737, A2 => n31144, B1 => n31141, B2 => 
                           n31133, ZN => n7880);
   U23619 : OAI22_X1 port map( A1 => n30855, A2 => n25526, B1 => n31125, B2 => 
                           n30848, ZN => n7365);
   U23620 : OAI22_X1 port map( A1 => n30855, A2 => n25525, B1 => n31128, B2 => 
                           n30848, ZN => n7366);
   U23621 : OAI22_X1 port map( A1 => n30855, A2 => n25524, B1 => n31131, B2 => 
                           n30848, ZN => n7367);
   U23622 : OAI22_X1 port map( A1 => n30855, A2 => n25522, B1 => n31134, B2 => 
                           n30848, ZN => n7368);
   U23623 : OAI22_X1 port map( A1 => n17776, A2 => n30779, B1 => n31125, B2 => 
                           n30773, ZN => n6981);
   U23624 : OAI22_X1 port map( A1 => n17775, A2 => n30779, B1 => n31128, B2 => 
                           n30773, ZN => n6982);
   U23625 : OAI22_X1 port map( A1 => n17774, A2 => n30779, B1 => n31131, B2 => 
                           n30773, ZN => n6983);
   U23626 : OAI22_X1 port map( A1 => n17772, A2 => n30779, B1 => n31134, B2 => 
                           n30773, ZN => n6984);
   U23627 : OAI22_X1 port map( A1 => n30931, A2 => n25241, B1 => n31124, B2 => 
                           n30924, ZN => n7749);
   U23628 : OAI22_X1 port map( A1 => n30931, A2 => n25240, B1 => n31127, B2 => 
                           n30924, ZN => n7750);
   U23629 : OAI22_X1 port map( A1 => n30931, A2 => n25239, B1 => n31130, B2 => 
                           n30924, ZN => n7751);
   U23630 : OAI22_X1 port map( A1 => n30931, A2 => n25237, B1 => n31133, B2 => 
                           n30924, ZN => n7752);
   U23631 : OAI22_X1 port map( A1 => n30881, A2 => n25390, B1 => n31124, B2 => 
                           n30874, ZN => n7493);
   U23632 : OAI22_X1 port map( A1 => n30881, A2 => n25389, B1 => n31127, B2 => 
                           n30874, ZN => n7494);
   U23633 : OAI22_X1 port map( A1 => n30881, A2 => n25388, B1 => n31130, B2 => 
                           n30874, ZN => n7495);
   U23634 : OAI22_X1 port map( A1 => n30881, A2 => n25386, B1 => n31133, B2 => 
                           n30874, ZN => n7496);
   U23635 : OAI22_X1 port map( A1 => n18063, A2 => n30679, B1 => n31125, B2 => 
                           n30673, ZN => n6469);
   U23636 : OAI22_X1 port map( A1 => n18062, A2 => n30679, B1 => n31128, B2 => 
                           n30673, ZN => n6470);
   U23637 : OAI22_X1 port map( A1 => n18061, A2 => n30679, B1 => n31131, B2 => 
                           n30673, ZN => n6471);
   U23638 : OAI22_X1 port map( A1 => n18059, A2 => n30679, B1 => n31134, B2 => 
                           n30673, ZN => n6472);
   U23639 : OAI22_X1 port map( A1 => n30755, A2 => n25812, B1 => n31125, B2 => 
                           n30748, ZN => n6853);
   U23640 : OAI22_X1 port map( A1 => n30755, A2 => n25811, B1 => n31128, B2 => 
                           n30748, ZN => n6854);
   U23641 : OAI22_X1 port map( A1 => n30755, A2 => n25810, B1 => n31131, B2 => 
                           n30748, ZN => n6855);
   U23642 : OAI22_X1 port map( A1 => n30755, A2 => n25808, B1 => n31134, B2 => 
                           n30748, ZN => n6856);
   U23643 : OAI22_X1 port map( A1 => n18263, A2 => n30643, B1 => n31126, B2 => 
                           n30637, ZN => n6277);
   U23644 : OAI22_X1 port map( A1 => n18262, A2 => n30643, B1 => n31129, B2 => 
                           n30637, ZN => n6278);
   U23645 : OAI22_X1 port map( A1 => n18261, A2 => n30643, B1 => n31132, B2 => 
                           n30637, ZN => n6279);
   U23646 : OAI22_X1 port map( A1 => n18259, A2 => n30643, B1 => n31135, B2 => 
                           n30637, ZN => n6280);
   U23647 : OAI22_X1 port map( A1 => n18130, A2 => n30667, B1 => n31126, B2 => 
                           n30661, ZN => n6405);
   U23648 : OAI22_X1 port map( A1 => n18129, A2 => n30667, B1 => n31129, B2 => 
                           n30661, ZN => n6406);
   U23649 : OAI22_X1 port map( A1 => n18128, A2 => n30667, B1 => n31132, B2 => 
                           n30661, ZN => n6407);
   U23650 : OAI22_X1 port map( A1 => n18126, A2 => n30667, B1 => n31135, B2 => 
                           n30661, ZN => n6408);
   U23651 : OAI22_X1 port map( A1 => n30631, A2 => n26107, B1 => n31126, B2 => 
                           n30624, ZN => n6213);
   U23652 : OAI22_X1 port map( A1 => n30631, A2 => n26106, B1 => n31129, B2 => 
                           n30624, ZN => n6214);
   U23653 : OAI22_X1 port map( A1 => n30631, A2 => n26105, B1 => n31132, B2 => 
                           n30624, ZN => n6215);
   U23654 : OAI22_X1 port map( A1 => n30631, A2 => n26103, B1 => n31135, B2 => 
                           n30624, ZN => n6216);
   U23655 : OAI22_X1 port map( A1 => n18196, A2 => n30655, B1 => n31126, B2 => 
                           n30649, ZN => n6341);
   U23656 : OAI22_X1 port map( A1 => n18195, A2 => n30655, B1 => n31129, B2 => 
                           n30649, ZN => n6342);
   U23657 : OAI22_X1 port map( A1 => n18194, A2 => n30655, B1 => n31132, B2 => 
                           n30649, ZN => n6343);
   U23658 : OAI22_X1 port map( A1 => n18192, A2 => n30655, B1 => n31135, B2 => 
                           n30649, ZN => n6344);
   U23659 : OAI22_X1 port map( A1 => n8987, A2 => n30593, B1 => n31126, B2 => 
                           n30587, ZN => n6021);
   U23660 : OAI22_X1 port map( A1 => n8982, A2 => n30593, B1 => n31129, B2 => 
                           n30587, ZN => n6022);
   U23661 : OAI22_X1 port map( A1 => n8977, A2 => n30593, B1 => n31132, B2 => 
                           n30587, ZN => n6023);
   U23662 : OAI22_X1 port map( A1 => n8972, A2 => n30593, B1 => n31135, B2 => 
                           n30587, ZN => n6024);
   U23663 : OAI22_X1 port map( A1 => n9755, A2 => n30600, B1 => n31126, B2 => 
                           n30599, ZN => n6085);
   U23664 : OAI22_X1 port map( A1 => n9750, A2 => n30600, B1 => n31129, B2 => 
                           n30599, ZN => n6086);
   U23665 : OAI22_X1 port map( A1 => n9745, A2 => n30600, B1 => n31132, B2 => 
                           n30599, ZN => n6087);
   U23666 : OAI22_X1 port map( A1 => n9740, A2 => n30602, B1 => n31135, B2 => 
                           n30599, ZN => n6088);
   U23667 : OAI22_X1 port map( A1 => n30618, A2 => n26173, B1 => n31126, B2 => 
                           n30611, ZN => n6149);
   U23668 : OAI22_X1 port map( A1 => n30618, A2 => n26172, B1 => n31129, B2 => 
                           n30611, ZN => n6150);
   U23669 : OAI22_X1 port map( A1 => n30618, A2 => n26171, B1 => n31132, B2 => 
                           n30611, ZN => n6151);
   U23670 : OAI22_X1 port map( A1 => n30618, A2 => n26169, B1 => n31135, B2 => 
                           n30611, ZN => n6152);
   U23671 : OAI22_X1 port map( A1 => n8988, A2 => n30717, B1 => n31125, B2 => 
                           n30711, ZN => n6661);
   U23672 : OAI22_X1 port map( A1 => n8983, A2 => n30717, B1 => n31128, B2 => 
                           n30711, ZN => n6662);
   U23673 : OAI22_X1 port map( A1 => n8978, A2 => n30717, B1 => n31131, B2 => 
                           n30711, ZN => n6663);
   U23674 : OAI22_X1 port map( A1 => n8973, A2 => n30717, B1 => n31134, B2 => 
                           n30711, ZN => n6664);
   U23675 : OAI22_X1 port map( A1 => n9756, A2 => n30724, B1 => n31125, B2 => 
                           n30723, ZN => n6725);
   U23676 : OAI22_X1 port map( A1 => n9751, A2 => n30724, B1 => n31128, B2 => 
                           n30723, ZN => n6726);
   U23677 : OAI22_X1 port map( A1 => n9746, A2 => n30724, B1 => n31131, B2 => 
                           n30723, ZN => n6727);
   U23678 : OAI22_X1 port map( A1 => n9741, A2 => n30726, B1 => n31134, B2 => 
                           n30723, ZN => n6728);
   U23679 : OAI22_X1 port map( A1 => n30742, A2 => n25879, B1 => n31125, B2 => 
                           n30735, ZN => n6789);
   U23680 : OAI22_X1 port map( A1 => n30742, A2 => n25878, B1 => n31128, B2 => 
                           n30735, ZN => n6790);
   U23681 : OAI22_X1 port map( A1 => n30742, A2 => n25877, B1 => n31131, B2 => 
                           n30735, ZN => n6791);
   U23682 : OAI22_X1 port map( A1 => n30742, A2 => n25875, B1 => n31134, B2 => 
                           n30735, ZN => n6792);
   U23683 : OAI22_X1 port map( A1 => n9612, A2 => n30767, B1 => n31125, B2 => 
                           n30761, ZN => n6917);
   U23684 : OAI22_X1 port map( A1 => n9611, A2 => n30767, B1 => n31128, B2 => 
                           n30761, ZN => n6918);
   U23685 : OAI22_X1 port map( A1 => n9610, A2 => n30767, B1 => n31131, B2 => 
                           n30761, ZN => n6919);
   U23686 : OAI22_X1 port map( A1 => n9609, A2 => n30767, B1 => n31134, B2 => 
                           n30761, ZN => n6920);
   U23687 : OAI22_X1 port map( A1 => n8986, A2 => n30817, B1 => n31125, B2 => 
                           n30811, ZN => n7173);
   U23688 : OAI22_X1 port map( A1 => n8981, A2 => n30817, B1 => n31128, B2 => 
                           n30811, ZN => n7174);
   U23689 : OAI22_X1 port map( A1 => n8976, A2 => n30817, B1 => n31131, B2 => 
                           n30811, ZN => n7175);
   U23690 : OAI22_X1 port map( A1 => n8971, A2 => n30817, B1 => n31134, B2 => 
                           n30811, ZN => n7176);
   U23691 : OAI22_X1 port map( A1 => n9754, A2 => n30824, B1 => n31124, B2 => 
                           n30823, ZN => n7237);
   U23692 : OAI22_X1 port map( A1 => n9749, A2 => n30824, B1 => n31127, B2 => 
                           n30823, ZN => n7238);
   U23693 : OAI22_X1 port map( A1 => n9744, A2 => n30824, B1 => n31130, B2 => 
                           n30823, ZN => n7239);
   U23694 : OAI22_X1 port map( A1 => n9739, A2 => n30826, B1 => n31133, B2 => 
                           n30823, ZN => n7240);
   U23695 : OAI22_X1 port map( A1 => n30842, A2 => n25593, B1 => n31124, B2 => 
                           n30835, ZN => n7301);
   U23696 : OAI22_X1 port map( A1 => n30842, A2 => n25592, B1 => n31127, B2 => 
                           n30835, ZN => n7302);
   U23697 : OAI22_X1 port map( A1 => n30842, A2 => n25591, B1 => n31130, B2 => 
                           n30835, ZN => n7303);
   U23698 : OAI22_X1 port map( A1 => n30842, A2 => n25589, B1 => n31133, B2 => 
                           n30835, ZN => n7304);
   U23699 : OAI22_X1 port map( A1 => n30868, A2 => n25460, B1 => n31124, B2 => 
                           n30861, ZN => n7429);
   U23700 : OAI22_X1 port map( A1 => n30868, A2 => n25459, B1 => n31127, B2 => 
                           n30861, ZN => n7430);
   U23701 : OAI22_X1 port map( A1 => n30868, A2 => n25458, B1 => n31130, B2 => 
                           n30861, ZN => n7431);
   U23702 : OAI22_X1 port map( A1 => n30868, A2 => n25456, B1 => n31133, B2 => 
                           n30861, ZN => n7432);
   U23703 : OAI22_X1 port map( A1 => n8985, A2 => n30893, B1 => n31124, B2 => 
                           n30887, ZN => n7557);
   U23704 : OAI22_X1 port map( A1 => n8980, A2 => n30893, B1 => n31127, B2 => 
                           n30887, ZN => n7558);
   U23705 : OAI22_X1 port map( A1 => n8975, A2 => n30893, B1 => n31130, B2 => 
                           n30887, ZN => n7559);
   U23706 : OAI22_X1 port map( A1 => n8970, A2 => n30893, B1 => n31133, B2 => 
                           n30887, ZN => n7560);
   U23707 : OAI22_X1 port map( A1 => n9753, A2 => n30900, B1 => n31124, B2 => 
                           n30899, ZN => n7621);
   U23708 : OAI22_X1 port map( A1 => n9748, A2 => n30900, B1 => n31127, B2 => 
                           n30899, ZN => n7622);
   U23709 : OAI22_X1 port map( A1 => n9743, A2 => n30900, B1 => n31130, B2 => 
                           n30899, ZN => n7623);
   U23710 : OAI22_X1 port map( A1 => n9738, A2 => n30902, B1 => n31133, B2 => 
                           n30899, ZN => n7624);
   U23711 : OAI22_X1 port map( A1 => n30918, A2 => n25308, B1 => n31124, B2 => 
                           n30911, ZN => n7685);
   U23712 : OAI22_X1 port map( A1 => n30918, A2 => n25307, B1 => n31127, B2 => 
                           n30911, ZN => n7686);
   U23713 : OAI22_X1 port map( A1 => n30918, A2 => n25306, B1 => n31130, B2 => 
                           n30911, ZN => n7687);
   U23714 : OAI22_X1 port map( A1 => n30918, A2 => n25304, B1 => n31133, B2 => 
                           n30911, ZN => n7688);
   U23715 : OAI22_X1 port map( A1 => n8984, A2 => n30943, B1 => n31124, B2 => 
                           n30937, ZN => n7813);
   U23716 : OAI22_X1 port map( A1 => n8979, A2 => n30943, B1 => n31127, B2 => 
                           n30937, ZN => n7814);
   U23717 : OAI22_X1 port map( A1 => n8974, A2 => n30943, B1 => n31130, B2 => 
                           n30937, ZN => n7815);
   U23718 : OAI22_X1 port map( A1 => n8969, A2 => n30943, B1 => n31133, B2 => 
                           n30937, ZN => n7816);
   U23719 : INV_X1 port map( A => ADD_RD1(4), ZN => n29306);
   U23720 : INV_X1 port map( A => ADD_RD2(4), ZN => n28029);
   U23721 : OAI22_X1 port map( A1 => n18244, A2 => n30651, B1 => n30982, B2 => 
                           n30645, ZN => n6293);
   U23722 : OAI22_X1 port map( A1 => n18243, A2 => n30651, B1 => n30985, B2 => 
                           n30645, ZN => n6294);
   U23723 : OAI22_X1 port map( A1 => n18242, A2 => n30651, B1 => n30988, B2 => 
                           n30645, ZN => n6295);
   U23724 : OAI22_X1 port map( A1 => n18241, A2 => n30651, B1 => n30991, B2 => 
                           n30645, ZN => n6296);
   U23725 : OAI22_X1 port map( A1 => n18240, A2 => n30651, B1 => n30994, B2 => 
                           n30645, ZN => n6297);
   U23726 : OAI22_X1 port map( A1 => n18239, A2 => n30651, B1 => n30997, B2 => 
                           n30645, ZN => n6298);
   U23727 : OAI22_X1 port map( A1 => n18238, A2 => n30651, B1 => n31000, B2 => 
                           n30645, ZN => n6299);
   U23728 : OAI22_X1 port map( A1 => n18237, A2 => n30651, B1 => n31003, B2 => 
                           n30645, ZN => n6300);
   U23729 : OAI22_X1 port map( A1 => n18236, A2 => n30651, B1 => n31006, B2 => 
                           n30645, ZN => n6301);
   U23730 : OAI22_X1 port map( A1 => n18235, A2 => n30651, B1 => n31009, B2 => 
                           n30645, ZN => n6302);
   U23731 : OAI22_X1 port map( A1 => n18234, A2 => n30651, B1 => n31012, B2 => 
                           n30645, ZN => n6303);
   U23732 : OAI22_X1 port map( A1 => n18233, A2 => n30652, B1 => n31015, B2 => 
                           n30645, ZN => n6304);
   U23733 : OAI22_X1 port map( A1 => n18232, A2 => n30652, B1 => n31018, B2 => 
                           n30646, ZN => n6305);
   U23734 : OAI22_X1 port map( A1 => n18231, A2 => n30652, B1 => n31021, B2 => 
                           n30646, ZN => n6306);
   U23735 : OAI22_X1 port map( A1 => n18230, A2 => n30652, B1 => n31024, B2 => 
                           n30646, ZN => n6307);
   U23736 : OAI22_X1 port map( A1 => n18229, A2 => n30652, B1 => n31027, B2 => 
                           n30646, ZN => n6308);
   U23737 : OAI22_X1 port map( A1 => n18228, A2 => n30652, B1 => n31030, B2 => 
                           n30646, ZN => n6309);
   U23738 : OAI22_X1 port map( A1 => n18227, A2 => n30652, B1 => n31033, B2 => 
                           n30646, ZN => n6310);
   U23739 : OAI22_X1 port map( A1 => n18226, A2 => n30652, B1 => n31036, B2 => 
                           n30646, ZN => n6311);
   U23740 : OAI22_X1 port map( A1 => n18225, A2 => n30652, B1 => n31039, B2 => 
                           n30646, ZN => n6312);
   U23741 : OAI22_X1 port map( A1 => n18224, A2 => n30652, B1 => n31042, B2 => 
                           n30646, ZN => n6313);
   U23742 : OAI22_X1 port map( A1 => n18223, A2 => n30652, B1 => n31045, B2 => 
                           n30646, ZN => n6314);
   U23743 : OAI22_X1 port map( A1 => n18222, A2 => n30652, B1 => n31048, B2 => 
                           n30646, ZN => n6315);
   U23744 : OAI22_X1 port map( A1 => n18221, A2 => n30653, B1 => n31051, B2 => 
                           n30646, ZN => n6316);
   U23745 : OAI22_X1 port map( A1 => n18220, A2 => n30653, B1 => n31054, B2 => 
                           n30647, ZN => n6317);
   U23746 : OAI22_X1 port map( A1 => n18219, A2 => n30653, B1 => n31057, B2 => 
                           n30647, ZN => n6318);
   U23747 : OAI22_X1 port map( A1 => n18311, A2 => n30639, B1 => n30982, B2 => 
                           n30633, ZN => n6229);
   U23748 : OAI22_X1 port map( A1 => n18310, A2 => n30639, B1 => n30985, B2 => 
                           n30633, ZN => n6230);
   U23749 : OAI22_X1 port map( A1 => n18309, A2 => n30639, B1 => n30988, B2 => 
                           n30633, ZN => n6231);
   U23750 : OAI22_X1 port map( A1 => n18308, A2 => n30639, B1 => n30991, B2 => 
                           n30633, ZN => n6232);
   U23751 : OAI22_X1 port map( A1 => n18307, A2 => n30639, B1 => n30994, B2 => 
                           n30633, ZN => n6233);
   U23752 : OAI22_X1 port map( A1 => n18306, A2 => n30639, B1 => n30997, B2 => 
                           n30633, ZN => n6234);
   U23753 : OAI22_X1 port map( A1 => n18305, A2 => n30639, B1 => n31000, B2 => 
                           n30633, ZN => n6235);
   U23754 : OAI22_X1 port map( A1 => n18304, A2 => n30639, B1 => n31003, B2 => 
                           n30633, ZN => n6236);
   U23755 : OAI22_X1 port map( A1 => n18303, A2 => n30639, B1 => n31006, B2 => 
                           n30633, ZN => n6237);
   U23756 : OAI22_X1 port map( A1 => n18302, A2 => n30639, B1 => n31009, B2 => 
                           n30633, ZN => n6238);
   U23757 : OAI22_X1 port map( A1 => n18301, A2 => n30639, B1 => n31012, B2 => 
                           n30633, ZN => n6239);
   U23758 : OAI22_X1 port map( A1 => n18300, A2 => n30640, B1 => n31015, B2 => 
                           n30633, ZN => n6240);
   U23759 : OAI22_X1 port map( A1 => n18299, A2 => n30640, B1 => n31018, B2 => 
                           n30634, ZN => n6241);
   U23760 : OAI22_X1 port map( A1 => n18298, A2 => n30640, B1 => n31021, B2 => 
                           n30634, ZN => n6242);
   U23761 : OAI22_X1 port map( A1 => n18297, A2 => n30640, B1 => n31024, B2 => 
                           n30634, ZN => n6243);
   U23762 : OAI22_X1 port map( A1 => n18296, A2 => n30640, B1 => n31027, B2 => 
                           n30634, ZN => n6244);
   U23763 : OAI22_X1 port map( A1 => n18295, A2 => n30640, B1 => n31030, B2 => 
                           n30634, ZN => n6245);
   U23764 : OAI22_X1 port map( A1 => n18294, A2 => n30640, B1 => n31033, B2 => 
                           n30634, ZN => n6246);
   U23765 : OAI22_X1 port map( A1 => n18293, A2 => n30640, B1 => n31036, B2 => 
                           n30634, ZN => n6247);
   U23766 : OAI22_X1 port map( A1 => n18292, A2 => n30640, B1 => n31039, B2 => 
                           n30634, ZN => n6248);
   U23767 : OAI22_X1 port map( A1 => n18291, A2 => n30640, B1 => n31042, B2 => 
                           n30634, ZN => n6249);
   U23768 : OAI22_X1 port map( A1 => n18290, A2 => n30640, B1 => n31045, B2 => 
                           n30634, ZN => n6250);
   U23769 : OAI22_X1 port map( A1 => n18289, A2 => n30640, B1 => n31048, B2 => 
                           n30634, ZN => n6251);
   U23770 : OAI22_X1 port map( A1 => n18288, A2 => n30641, B1 => n31051, B2 => 
                           n30634, ZN => n6252);
   U23771 : OAI22_X1 port map( A1 => n18287, A2 => n30641, B1 => n31054, B2 => 
                           n30635, ZN => n6253);
   U23772 : OAI22_X1 port map( A1 => n18286, A2 => n30641, B1 => n31057, B2 => 
                           n30635, ZN => n6254);
   U23773 : OAI22_X1 port map( A1 => n18218, A2 => n30653, B1 => n31060, B2 => 
                           n30647, ZN => n6319);
   U23774 : OAI22_X1 port map( A1 => n18217, A2 => n30653, B1 => n31063, B2 => 
                           n30647, ZN => n6320);
   U23775 : OAI22_X1 port map( A1 => n18216, A2 => n30653, B1 => n31066, B2 => 
                           n30647, ZN => n6321);
   U23776 : OAI22_X1 port map( A1 => n18215, A2 => n30653, B1 => n31069, B2 => 
                           n30647, ZN => n6322);
   U23777 : OAI22_X1 port map( A1 => n18214, A2 => n30653, B1 => n31072, B2 => 
                           n30647, ZN => n6323);
   U23778 : OAI22_X1 port map( A1 => n18213, A2 => n30653, B1 => n31075, B2 => 
                           n30647, ZN => n6324);
   U23779 : OAI22_X1 port map( A1 => n18212, A2 => n30653, B1 => n31078, B2 => 
                           n30647, ZN => n6325);
   U23780 : OAI22_X1 port map( A1 => n18211, A2 => n30653, B1 => n31081, B2 => 
                           n30647, ZN => n6326);
   U23781 : OAI22_X1 port map( A1 => n18210, A2 => n30653, B1 => n31084, B2 => 
                           n30647, ZN => n6327);
   U23782 : OAI22_X1 port map( A1 => n18209, A2 => n30654, B1 => n31087, B2 => 
                           n30647, ZN => n6328);
   U23783 : OAI22_X1 port map( A1 => n18208, A2 => n30654, B1 => n31090, B2 => 
                           n30648, ZN => n6329);
   U23784 : OAI22_X1 port map( A1 => n18207, A2 => n30654, B1 => n31093, B2 => 
                           n30648, ZN => n6330);
   U23785 : OAI22_X1 port map( A1 => n18206, A2 => n30654, B1 => n31096, B2 => 
                           n30648, ZN => n6331);
   U23786 : OAI22_X1 port map( A1 => n18205, A2 => n30654, B1 => n31099, B2 => 
                           n30648, ZN => n6332);
   U23787 : OAI22_X1 port map( A1 => n18204, A2 => n30654, B1 => n31102, B2 => 
                           n30648, ZN => n6333);
   U23788 : OAI22_X1 port map( A1 => n18203, A2 => n30654, B1 => n31105, B2 => 
                           n30648, ZN => n6334);
   U23789 : OAI22_X1 port map( A1 => n18202, A2 => n30654, B1 => n31108, B2 => 
                           n30648, ZN => n6335);
   U23790 : OAI22_X1 port map( A1 => n18201, A2 => n30654, B1 => n31111, B2 => 
                           n30648, ZN => n6336);
   U23791 : OAI22_X1 port map( A1 => n18200, A2 => n30654, B1 => n31114, B2 => 
                           n30648, ZN => n6337);
   U23792 : OAI22_X1 port map( A1 => n18199, A2 => n30654, B1 => n31117, B2 => 
                           n30648, ZN => n6338);
   U23793 : OAI22_X1 port map( A1 => n18198, A2 => n30654, B1 => n31120, B2 => 
                           n30648, ZN => n6339);
   U23794 : OAI22_X1 port map( A1 => n18197, A2 => n30655, B1 => n31123, B2 => 
                           n30648, ZN => n6340);
   U23795 : OAI22_X1 port map( A1 => n18285, A2 => n30641, B1 => n31060, B2 => 
                           n30635, ZN => n6255);
   U23796 : OAI22_X1 port map( A1 => n18284, A2 => n30641, B1 => n31063, B2 => 
                           n30635, ZN => n6256);
   U23797 : OAI22_X1 port map( A1 => n18283, A2 => n30641, B1 => n31066, B2 => 
                           n30635, ZN => n6257);
   U23798 : OAI22_X1 port map( A1 => n18282, A2 => n30641, B1 => n31069, B2 => 
                           n30635, ZN => n6258);
   U23799 : OAI22_X1 port map( A1 => n18281, A2 => n30641, B1 => n31072, B2 => 
                           n30635, ZN => n6259);
   U23800 : OAI22_X1 port map( A1 => n18280, A2 => n30641, B1 => n31075, B2 => 
                           n30635, ZN => n6260);
   U23801 : OAI22_X1 port map( A1 => n18279, A2 => n30641, B1 => n31078, B2 => 
                           n30635, ZN => n6261);
   U23802 : OAI22_X1 port map( A1 => n18278, A2 => n30641, B1 => n31081, B2 => 
                           n30635, ZN => n6262);
   U23803 : OAI22_X1 port map( A1 => n18277, A2 => n30641, B1 => n31084, B2 => 
                           n30635, ZN => n6263);
   U23804 : OAI22_X1 port map( A1 => n18276, A2 => n30642, B1 => n31087, B2 => 
                           n30635, ZN => n6264);
   U23805 : OAI22_X1 port map( A1 => n18275, A2 => n30642, B1 => n31090, B2 => 
                           n30636, ZN => n6265);
   U23806 : OAI22_X1 port map( A1 => n18274, A2 => n30642, B1 => n31093, B2 => 
                           n30636, ZN => n6266);
   U23807 : OAI22_X1 port map( A1 => n18273, A2 => n30642, B1 => n31096, B2 => 
                           n30636, ZN => n6267);
   U23808 : OAI22_X1 port map( A1 => n18272, A2 => n30642, B1 => n31099, B2 => 
                           n30636, ZN => n6268);
   U23809 : OAI22_X1 port map( A1 => n18271, A2 => n30642, B1 => n31102, B2 => 
                           n30636, ZN => n6269);
   U23810 : OAI22_X1 port map( A1 => n18270, A2 => n30642, B1 => n31105, B2 => 
                           n30636, ZN => n6270);
   U23811 : OAI22_X1 port map( A1 => n18269, A2 => n30642, B1 => n31108, B2 => 
                           n30636, ZN => n6271);
   U23812 : OAI22_X1 port map( A1 => n18268, A2 => n30642, B1 => n31111, B2 => 
                           n30636, ZN => n6272);
   U23813 : OAI22_X1 port map( A1 => n18267, A2 => n30642, B1 => n31114, B2 => 
                           n30636, ZN => n6273);
   U23814 : OAI22_X1 port map( A1 => n18266, A2 => n30642, B1 => n31117, B2 => 
                           n30636, ZN => n6274);
   U23815 : OAI22_X1 port map( A1 => n18265, A2 => n30642, B1 => n31120, B2 => 
                           n30636, ZN => n6275);
   U23816 : OAI22_X1 port map( A1 => n18264, A2 => n30643, B1 => n31123, B2 => 
                           n30636, ZN => n6276);
   U23817 : OAI22_X1 port map( A1 => n18256, A2 => n30650, B1 => n30946, B2 => 
                           n30644, ZN => n6281);
   U23818 : OAI22_X1 port map( A1 => n18255, A2 => n30650, B1 => n30949, B2 => 
                           n30644, ZN => n6282);
   U23819 : OAI22_X1 port map( A1 => n18254, A2 => n30650, B1 => n30952, B2 => 
                           n30644, ZN => n6283);
   U23820 : OAI22_X1 port map( A1 => n18253, A2 => n30650, B1 => n30955, B2 => 
                           n30644, ZN => n6284);
   U23821 : OAI22_X1 port map( A1 => n18252, A2 => n30650, B1 => n30958, B2 => 
                           n30644, ZN => n6285);
   U23822 : OAI22_X1 port map( A1 => n18251, A2 => n30650, B1 => n30961, B2 => 
                           n30644, ZN => n6286);
   U23823 : OAI22_X1 port map( A1 => n18250, A2 => n30650, B1 => n30964, B2 => 
                           n30644, ZN => n6287);
   U23824 : OAI22_X1 port map( A1 => n18249, A2 => n30650, B1 => n30967, B2 => 
                           n30644, ZN => n6288);
   U23825 : OAI22_X1 port map( A1 => n18248, A2 => n30650, B1 => n30970, B2 => 
                           n30644, ZN => n6289);
   U23826 : OAI22_X1 port map( A1 => n18247, A2 => n30650, B1 => n30973, B2 => 
                           n30644, ZN => n6290);
   U23827 : OAI22_X1 port map( A1 => n18246, A2 => n30650, B1 => n30976, B2 => 
                           n30644, ZN => n6291);
   U23828 : OAI22_X1 port map( A1 => n18245, A2 => n30651, B1 => n30979, B2 => 
                           n30644, ZN => n6292);
   U23829 : OAI22_X1 port map( A1 => n18323, A2 => n30638, B1 => n30946, B2 => 
                           n30632, ZN => n6217);
   U23830 : OAI22_X1 port map( A1 => n18322, A2 => n30638, B1 => n30949, B2 => 
                           n30632, ZN => n6218);
   U23831 : OAI22_X1 port map( A1 => n18321, A2 => n30638, B1 => n30952, B2 => 
                           n30632, ZN => n6219);
   U23832 : OAI22_X1 port map( A1 => n18320, A2 => n30638, B1 => n30955, B2 => 
                           n30632, ZN => n6220);
   U23833 : OAI22_X1 port map( A1 => n18319, A2 => n30638, B1 => n30958, B2 => 
                           n30632, ZN => n6221);
   U23834 : OAI22_X1 port map( A1 => n18318, A2 => n30638, B1 => n30961, B2 => 
                           n30632, ZN => n6222);
   U23835 : OAI22_X1 port map( A1 => n18317, A2 => n30638, B1 => n30964, B2 => 
                           n30632, ZN => n6223);
   U23836 : OAI22_X1 port map( A1 => n18316, A2 => n30638, B1 => n30967, B2 => 
                           n30632, ZN => n6224);
   U23837 : OAI22_X1 port map( A1 => n18315, A2 => n30638, B1 => n30970, B2 => 
                           n30632, ZN => n6225);
   U23838 : OAI22_X1 port map( A1 => n18314, A2 => n30638, B1 => n30973, B2 => 
                           n30632, ZN => n6226);
   U23839 : OAI22_X1 port map( A1 => n18313, A2 => n30638, B1 => n30976, B2 => 
                           n30632, ZN => n6227);
   U23840 : OAI22_X1 port map( A1 => n18312, A2 => n30639, B1 => n30979, B2 => 
                           n30632, ZN => n6228);
   U23841 : OAI22_X1 port map( A1 => n30628, A2 => n26155, B1 => n30982, B2 => 
                           n30620, ZN => n6165);
   U23842 : OAI22_X1 port map( A1 => n30628, A2 => n26154, B1 => n30985, B2 => 
                           n30620, ZN => n6166);
   U23843 : OAI22_X1 port map( A1 => n30628, A2 => n26153, B1 => n30988, B2 => 
                           n30620, ZN => n6167);
   U23844 : OAI22_X1 port map( A1 => n30628, A2 => n26152, B1 => n30991, B2 => 
                           n30620, ZN => n6168);
   U23845 : OAI22_X1 port map( A1 => n30628, A2 => n26151, B1 => n30994, B2 => 
                           n30620, ZN => n6169);
   U23846 : OAI22_X1 port map( A1 => n30628, A2 => n26150, B1 => n30997, B2 => 
                           n30620, ZN => n6170);
   U23847 : OAI22_X1 port map( A1 => n30628, A2 => n26149, B1 => n31000, B2 => 
                           n30620, ZN => n6171);
   U23848 : OAI22_X1 port map( A1 => n30628, A2 => n26148, B1 => n31003, B2 => 
                           n30620, ZN => n6172);
   U23849 : OAI22_X1 port map( A1 => n30628, A2 => n26147, B1 => n31006, B2 => 
                           n30620, ZN => n6173);
   U23850 : OAI22_X1 port map( A1 => n30628, A2 => n26146, B1 => n31009, B2 => 
                           n30620, ZN => n6174);
   U23851 : OAI22_X1 port map( A1 => n30628, A2 => n26145, B1 => n31012, B2 => 
                           n30620, ZN => n6175);
   U23852 : OAI22_X1 port map( A1 => n30628, A2 => n26144, B1 => n31015, B2 => 
                           n30620, ZN => n6176);
   U23853 : OAI22_X1 port map( A1 => n30628, A2 => n26143, B1 => n31018, B2 => 
                           n30621, ZN => n6177);
   U23854 : OAI22_X1 port map( A1 => n30629, A2 => n26142, B1 => n31021, B2 => 
                           n30621, ZN => n6178);
   U23855 : OAI22_X1 port map( A1 => n30629, A2 => n26141, B1 => n31024, B2 => 
                           n30621, ZN => n6179);
   U23856 : OAI22_X1 port map( A1 => n30629, A2 => n26140, B1 => n31027, B2 => 
                           n30621, ZN => n6180);
   U23857 : OAI22_X1 port map( A1 => n30629, A2 => n26139, B1 => n31030, B2 => 
                           n30621, ZN => n6181);
   U23858 : OAI22_X1 port map( A1 => n30629, A2 => n26138, B1 => n31033, B2 => 
                           n30621, ZN => n6182);
   U23859 : OAI22_X1 port map( A1 => n30629, A2 => n26137, B1 => n31036, B2 => 
                           n30621, ZN => n6183);
   U23860 : OAI22_X1 port map( A1 => n30629, A2 => n26136, B1 => n31039, B2 => 
                           n30621, ZN => n6184);
   U23861 : OAI22_X1 port map( A1 => n30629, A2 => n26135, B1 => n31042, B2 => 
                           n30621, ZN => n6185);
   U23862 : OAI22_X1 port map( A1 => n30629, A2 => n26134, B1 => n31045, B2 => 
                           n30621, ZN => n6186);
   U23863 : OAI22_X1 port map( A1 => n30629, A2 => n26133, B1 => n31048, B2 => 
                           n30621, ZN => n6187);
   U23864 : OAI22_X1 port map( A1 => n30629, A2 => n26132, B1 => n31051, B2 => 
                           n30621, ZN => n6188);
   U23865 : OAI22_X1 port map( A1 => n30629, A2 => n26131, B1 => n31054, B2 => 
                           n30622, ZN => n6189);
   U23866 : OAI22_X1 port map( A1 => n30629, A2 => n26130, B1 => n31057, B2 => 
                           n30622, ZN => n6190);
   U23867 : OAI22_X1 port map( A1 => n30630, A2 => n26129, B1 => n31060, B2 => 
                           n30622, ZN => n6191);
   U23868 : OAI22_X1 port map( A1 => n30630, A2 => n26128, B1 => n31063, B2 => 
                           n30622, ZN => n6192);
   U23869 : OAI22_X1 port map( A1 => n30630, A2 => n26127, B1 => n31066, B2 => 
                           n30622, ZN => n6193);
   U23870 : OAI22_X1 port map( A1 => n30630, A2 => n26126, B1 => n31069, B2 => 
                           n30622, ZN => n6194);
   U23871 : OAI22_X1 port map( A1 => n30630, A2 => n26125, B1 => n31072, B2 => 
                           n30622, ZN => n6195);
   U23872 : OAI22_X1 port map( A1 => n30630, A2 => n26124, B1 => n31075, B2 => 
                           n30622, ZN => n6196);
   U23873 : OAI22_X1 port map( A1 => n30630, A2 => n26123, B1 => n31078, B2 => 
                           n30622, ZN => n6197);
   U23874 : OAI22_X1 port map( A1 => n30630, A2 => n26122, B1 => n31081, B2 => 
                           n30622, ZN => n6198);
   U23875 : OAI22_X1 port map( A1 => n30630, A2 => n26121, B1 => n31084, B2 => 
                           n30622, ZN => n6199);
   U23876 : OAI22_X1 port map( A1 => n30630, A2 => n26120, B1 => n31087, B2 => 
                           n30622, ZN => n6200);
   U23877 : OAI22_X1 port map( A1 => n30630, A2 => n26119, B1 => n31090, B2 => 
                           n30623, ZN => n6201);
   U23878 : OAI22_X1 port map( A1 => n30630, A2 => n26118, B1 => n31093, B2 => 
                           n30623, ZN => n6202);
   U23879 : OAI22_X1 port map( A1 => n30630, A2 => n26117, B1 => n31096, B2 => 
                           n30623, ZN => n6203);
   U23880 : OAI22_X1 port map( A1 => n30631, A2 => n26116, B1 => n31099, B2 => 
                           n30623, ZN => n6204);
   U23881 : OAI22_X1 port map( A1 => n30631, A2 => n26115, B1 => n31102, B2 => 
                           n30623, ZN => n6205);
   U23882 : OAI22_X1 port map( A1 => n30631, A2 => n26114, B1 => n31105, B2 => 
                           n30623, ZN => n6206);
   U23883 : OAI22_X1 port map( A1 => n30631, A2 => n26113, B1 => n31108, B2 => 
                           n30623, ZN => n6207);
   U23884 : OAI22_X1 port map( A1 => n30631, A2 => n26112, B1 => n31111, B2 => 
                           n30623, ZN => n6208);
   U23885 : OAI22_X1 port map( A1 => n30631, A2 => n26111, B1 => n31114, B2 => 
                           n30623, ZN => n6209);
   U23886 : OAI22_X1 port map( A1 => n30631, A2 => n26110, B1 => n31117, B2 => 
                           n30623, ZN => n6210);
   U23887 : OAI22_X1 port map( A1 => n30631, A2 => n26109, B1 => n31120, B2 => 
                           n30623, ZN => n6211);
   U23888 : OAI22_X1 port map( A1 => n30631, A2 => n26108, B1 => n31123, B2 => 
                           n30623, ZN => n6212);
   U23889 : OAI22_X1 port map( A1 => n18178, A2 => n30663, B1 => n30982, B2 => 
                           n30657, ZN => n6357);
   U23890 : OAI22_X1 port map( A1 => n18177, A2 => n30663, B1 => n30985, B2 => 
                           n30657, ZN => n6358);
   U23891 : OAI22_X1 port map( A1 => n18176, A2 => n30663, B1 => n30988, B2 => 
                           n30657, ZN => n6359);
   U23892 : OAI22_X1 port map( A1 => n18175, A2 => n30663, B1 => n30991, B2 => 
                           n30657, ZN => n6360);
   U23893 : OAI22_X1 port map( A1 => n18174, A2 => n30663, B1 => n30994, B2 => 
                           n30657, ZN => n6361);
   U23894 : OAI22_X1 port map( A1 => n18173, A2 => n30663, B1 => n30997, B2 => 
                           n30657, ZN => n6362);
   U23895 : OAI22_X1 port map( A1 => n18172, A2 => n30663, B1 => n31000, B2 => 
                           n30657, ZN => n6363);
   U23896 : OAI22_X1 port map( A1 => n18171, A2 => n30663, B1 => n31003, B2 => 
                           n30657, ZN => n6364);
   U23897 : OAI22_X1 port map( A1 => n18170, A2 => n30663, B1 => n31006, B2 => 
                           n30657, ZN => n6365);
   U23898 : OAI22_X1 port map( A1 => n18169, A2 => n30663, B1 => n31009, B2 => 
                           n30657, ZN => n6366);
   U23899 : OAI22_X1 port map( A1 => n18168, A2 => n30663, B1 => n31012, B2 => 
                           n30657, ZN => n6367);
   U23900 : OAI22_X1 port map( A1 => n18167, A2 => n30664, B1 => n31015, B2 => 
                           n30657, ZN => n6368);
   U23901 : OAI22_X1 port map( A1 => n18166, A2 => n30664, B1 => n31018, B2 => 
                           n30658, ZN => n6369);
   U23902 : OAI22_X1 port map( A1 => n18165, A2 => n30664, B1 => n31021, B2 => 
                           n30658, ZN => n6370);
   U23903 : OAI22_X1 port map( A1 => n18164, A2 => n30664, B1 => n31024, B2 => 
                           n30658, ZN => n6371);
   U23904 : OAI22_X1 port map( A1 => n18163, A2 => n30664, B1 => n31027, B2 => 
                           n30658, ZN => n6372);
   U23905 : OAI22_X1 port map( A1 => n18162, A2 => n30664, B1 => n31030, B2 => 
                           n30658, ZN => n6373);
   U23906 : OAI22_X1 port map( A1 => n18161, A2 => n30664, B1 => n31033, B2 => 
                           n30658, ZN => n6374);
   U23907 : OAI22_X1 port map( A1 => n18160, A2 => n30664, B1 => n31036, B2 => 
                           n30658, ZN => n6375);
   U23908 : OAI22_X1 port map( A1 => n18159, A2 => n30664, B1 => n31039, B2 => 
                           n30658, ZN => n6376);
   U23909 : OAI22_X1 port map( A1 => n18158, A2 => n30664, B1 => n31042, B2 => 
                           n30658, ZN => n6377);
   U23910 : OAI22_X1 port map( A1 => n18157, A2 => n30664, B1 => n31045, B2 => 
                           n30658, ZN => n6378);
   U23911 : OAI22_X1 port map( A1 => n18156, A2 => n30664, B1 => n31048, B2 => 
                           n30658, ZN => n6379);
   U23912 : OAI22_X1 port map( A1 => n18155, A2 => n30665, B1 => n31051, B2 => 
                           n30658, ZN => n6380);
   U23913 : OAI22_X1 port map( A1 => n18154, A2 => n30665, B1 => n31054, B2 => 
                           n30659, ZN => n6381);
   U23914 : OAI22_X1 port map( A1 => n18153, A2 => n30665, B1 => n31057, B2 => 
                           n30659, ZN => n6382);
   U23915 : OAI22_X1 port map( A1 => n18152, A2 => n30665, B1 => n31060, B2 => 
                           n30659, ZN => n6383);
   U23916 : OAI22_X1 port map( A1 => n18151, A2 => n30665, B1 => n31063, B2 => 
                           n30659, ZN => n6384);
   U23917 : OAI22_X1 port map( A1 => n18150, A2 => n30665, B1 => n31066, B2 => 
                           n30659, ZN => n6385);
   U23918 : OAI22_X1 port map( A1 => n18149, A2 => n30665, B1 => n31069, B2 => 
                           n30659, ZN => n6386);
   U23919 : OAI22_X1 port map( A1 => n18148, A2 => n30665, B1 => n31072, B2 => 
                           n30659, ZN => n6387);
   U23920 : OAI22_X1 port map( A1 => n18147, A2 => n30665, B1 => n31075, B2 => 
                           n30659, ZN => n6388);
   U23921 : OAI22_X1 port map( A1 => n18146, A2 => n30665, B1 => n31078, B2 => 
                           n30659, ZN => n6389);
   U23922 : OAI22_X1 port map( A1 => n18145, A2 => n30665, B1 => n31081, B2 => 
                           n30659, ZN => n6390);
   U23923 : OAI22_X1 port map( A1 => n18144, A2 => n30665, B1 => n31084, B2 => 
                           n30659, ZN => n6391);
   U23924 : OAI22_X1 port map( A1 => n18143, A2 => n30666, B1 => n31087, B2 => 
                           n30659, ZN => n6392);
   U23925 : OAI22_X1 port map( A1 => n18142, A2 => n30666, B1 => n31090, B2 => 
                           n30660, ZN => n6393);
   U23926 : OAI22_X1 port map( A1 => n18141, A2 => n30666, B1 => n31093, B2 => 
                           n30660, ZN => n6394);
   U23927 : OAI22_X1 port map( A1 => n18140, A2 => n30666, B1 => n31096, B2 => 
                           n30660, ZN => n6395);
   U23928 : OAI22_X1 port map( A1 => n18139, A2 => n30666, B1 => n31099, B2 => 
                           n30660, ZN => n6396);
   U23929 : OAI22_X1 port map( A1 => n18138, A2 => n30666, B1 => n31102, B2 => 
                           n30660, ZN => n6397);
   U23930 : OAI22_X1 port map( A1 => n18137, A2 => n30666, B1 => n31105, B2 => 
                           n30660, ZN => n6398);
   U23931 : OAI22_X1 port map( A1 => n18136, A2 => n30666, B1 => n31108, B2 => 
                           n30660, ZN => n6399);
   U23932 : OAI22_X1 port map( A1 => n18135, A2 => n30666, B1 => n31111, B2 => 
                           n30660, ZN => n6400);
   U23933 : OAI22_X1 port map( A1 => n18134, A2 => n30666, B1 => n31114, B2 => 
                           n30660, ZN => n6401);
   U23934 : OAI22_X1 port map( A1 => n18133, A2 => n30666, B1 => n31117, B2 => 
                           n30660, ZN => n6402);
   U23935 : OAI22_X1 port map( A1 => n18132, A2 => n30666, B1 => n31120, B2 => 
                           n30660, ZN => n6403);
   U23936 : OAI22_X1 port map( A1 => n18131, A2 => n30667, B1 => n31123, B2 => 
                           n30660, ZN => n6404);
   U23937 : OAI22_X1 port map( A1 => n30627, A2 => n26167, B1 => n30946, B2 => 
                           n30619, ZN => n6153);
   U23938 : OAI22_X1 port map( A1 => n30627, A2 => n26166, B1 => n30949, B2 => 
                           n30619, ZN => n6154);
   U23939 : OAI22_X1 port map( A1 => n30627, A2 => n26165, B1 => n30952, B2 => 
                           n30619, ZN => n6155);
   U23940 : OAI22_X1 port map( A1 => n30627, A2 => n26164, B1 => n30955, B2 => 
                           n30619, ZN => n6156);
   U23941 : OAI22_X1 port map( A1 => n30627, A2 => n26163, B1 => n30958, B2 => 
                           n30619, ZN => n6157);
   U23942 : OAI22_X1 port map( A1 => n30627, A2 => n26162, B1 => n30961, B2 => 
                           n30619, ZN => n6158);
   U23943 : OAI22_X1 port map( A1 => n30627, A2 => n26161, B1 => n30964, B2 => 
                           n30619, ZN => n6159);
   U23944 : OAI22_X1 port map( A1 => n30627, A2 => n26160, B1 => n30967, B2 => 
                           n30619, ZN => n6160);
   U23945 : OAI22_X1 port map( A1 => n30627, A2 => n26159, B1 => n30970, B2 => 
                           n30619, ZN => n6161);
   U23946 : OAI22_X1 port map( A1 => n30627, A2 => n26158, B1 => n30973, B2 => 
                           n30619, ZN => n6162);
   U23947 : OAI22_X1 port map( A1 => n30627, A2 => n26157, B1 => n30976, B2 => 
                           n30619, ZN => n6163);
   U23948 : OAI22_X1 port map( A1 => n30627, A2 => n26156, B1 => n30979, B2 => 
                           n30619, ZN => n6164);
   U23949 : OAI22_X1 port map( A1 => n18190, A2 => n30662, B1 => n30946, B2 => 
                           n30656, ZN => n6345);
   U23950 : OAI22_X1 port map( A1 => n18189, A2 => n30662, B1 => n30949, B2 => 
                           n30656, ZN => n6346);
   U23951 : OAI22_X1 port map( A1 => n18188, A2 => n30662, B1 => n30952, B2 => 
                           n30656, ZN => n6347);
   U23952 : OAI22_X1 port map( A1 => n18187, A2 => n30662, B1 => n30955, B2 => 
                           n30656, ZN => n6348);
   U23953 : OAI22_X1 port map( A1 => n18186, A2 => n30662, B1 => n30958, B2 => 
                           n30656, ZN => n6349);
   U23954 : OAI22_X1 port map( A1 => n18185, A2 => n30662, B1 => n30961, B2 => 
                           n30656, ZN => n6350);
   U23955 : OAI22_X1 port map( A1 => n18184, A2 => n30662, B1 => n30964, B2 => 
                           n30656, ZN => n6351);
   U23956 : OAI22_X1 port map( A1 => n18183, A2 => n30662, B1 => n30967, B2 => 
                           n30656, ZN => n6352);
   U23957 : OAI22_X1 port map( A1 => n18182, A2 => n30662, B1 => n30970, B2 => 
                           n30656, ZN => n6353);
   U23958 : OAI22_X1 port map( A1 => n18181, A2 => n30662, B1 => n30973, B2 => 
                           n30656, ZN => n6354);
   U23959 : OAI22_X1 port map( A1 => n18180, A2 => n30662, B1 => n30976, B2 => 
                           n30656, ZN => n6355);
   U23960 : OAI22_X1 port map( A1 => n18179, A2 => n30663, B1 => n30979, B2 => 
                           n30656, ZN => n6356);
   U23961 : OAI22_X1 port map( A1 => n9287, A2 => n30588, B1 => n30946, B2 => 
                           n30582, ZN => n5961);
   U23962 : OAI22_X1 port map( A1 => n9282, A2 => n30588, B1 => n30949, B2 => 
                           n30582, ZN => n5962);
   U23963 : OAI22_X1 port map( A1 => n9277, A2 => n30588, B1 => n30952, B2 => 
                           n30582, ZN => n5963);
   U23964 : OAI22_X1 port map( A1 => n9272, A2 => n30588, B1 => n30955, B2 => 
                           n30582, ZN => n5964);
   U23965 : OAI22_X1 port map( A1 => n9267, A2 => n30588, B1 => n30958, B2 => 
                           n30582, ZN => n5965);
   U23966 : OAI22_X1 port map( A1 => n9262, A2 => n30588, B1 => n30961, B2 => 
                           n30582, ZN => n5966);
   U23967 : OAI22_X1 port map( A1 => n9257, A2 => n30588, B1 => n30964, B2 => 
                           n30582, ZN => n5967);
   U23968 : OAI22_X1 port map( A1 => n9252, A2 => n30588, B1 => n30967, B2 => 
                           n30582, ZN => n5968);
   U23969 : OAI22_X1 port map( A1 => n9247, A2 => n30588, B1 => n30970, B2 => 
                           n30582, ZN => n5969);
   U23970 : OAI22_X1 port map( A1 => n9242, A2 => n30588, B1 => n30973, B2 => 
                           n30582, ZN => n5970);
   U23971 : OAI22_X1 port map( A1 => n9237, A2 => n30588, B1 => n30976, B2 => 
                           n30582, ZN => n5971);
   U23972 : OAI22_X1 port map( A1 => n9232, A2 => n30589, B1 => n30979, B2 => 
                           n30582, ZN => n5972);
   U23973 : OAI22_X1 port map( A1 => n9227, A2 => n30589, B1 => n30982, B2 => 
                           n30583, ZN => n5973);
   U23974 : OAI22_X1 port map( A1 => n9222, A2 => n30589, B1 => n30985, B2 => 
                           n30583, ZN => n5974);
   U23975 : OAI22_X1 port map( A1 => n9217, A2 => n30589, B1 => n30988, B2 => 
                           n30583, ZN => n5975);
   U23976 : OAI22_X1 port map( A1 => n9212, A2 => n30589, B1 => n30991, B2 => 
                           n30583, ZN => n5976);
   U23977 : OAI22_X1 port map( A1 => n9207, A2 => n30589, B1 => n30994, B2 => 
                           n30583, ZN => n5977);
   U23978 : OAI22_X1 port map( A1 => n9202, A2 => n30589, B1 => n30997, B2 => 
                           n30583, ZN => n5978);
   U23979 : OAI22_X1 port map( A1 => n9197, A2 => n30589, B1 => n31000, B2 => 
                           n30583, ZN => n5979);
   U23980 : OAI22_X1 port map( A1 => n9192, A2 => n30589, B1 => n31003, B2 => 
                           n30583, ZN => n5980);
   U23981 : OAI22_X1 port map( A1 => n9187, A2 => n30589, B1 => n31006, B2 => 
                           n30583, ZN => n5981);
   U23982 : OAI22_X1 port map( A1 => n9182, A2 => n30589, B1 => n31009, B2 => 
                           n30583, ZN => n5982);
   U23983 : OAI22_X1 port map( A1 => n9177, A2 => n30589, B1 => n31012, B2 => 
                           n30583, ZN => n5983);
   U23984 : OAI22_X1 port map( A1 => n9172, A2 => n30590, B1 => n31015, B2 => 
                           n30583, ZN => n5984);
   U23985 : OAI22_X1 port map( A1 => n9167, A2 => n30590, B1 => n31018, B2 => 
                           n30584, ZN => n5985);
   U23986 : OAI22_X1 port map( A1 => n9162, A2 => n30590, B1 => n31021, B2 => 
                           n30584, ZN => n5986);
   U23987 : OAI22_X1 port map( A1 => n9157, A2 => n30590, B1 => n31024, B2 => 
                           n30584, ZN => n5987);
   U23988 : OAI22_X1 port map( A1 => n9152, A2 => n30590, B1 => n31027, B2 => 
                           n30584, ZN => n5988);
   U23989 : OAI22_X1 port map( A1 => n9147, A2 => n30590, B1 => n31030, B2 => 
                           n30584, ZN => n5989);
   U23990 : OAI22_X1 port map( A1 => n9142, A2 => n30590, B1 => n31033, B2 => 
                           n30584, ZN => n5990);
   U23991 : OAI22_X1 port map( A1 => n9137, A2 => n30590, B1 => n31036, B2 => 
                           n30584, ZN => n5991);
   U23992 : OAI22_X1 port map( A1 => n9132, A2 => n30590, B1 => n31039, B2 => 
                           n30584, ZN => n5992);
   U23993 : OAI22_X1 port map( A1 => n9127, A2 => n30590, B1 => n31042, B2 => 
                           n30584, ZN => n5993);
   U23994 : OAI22_X1 port map( A1 => n9122, A2 => n30590, B1 => n31045, B2 => 
                           n30584, ZN => n5994);
   U23995 : OAI22_X1 port map( A1 => n9117, A2 => n30590, B1 => n31048, B2 => 
                           n30584, ZN => n5995);
   U23996 : OAI22_X1 port map( A1 => n9112, A2 => n30591, B1 => n31051, B2 => 
                           n30584, ZN => n5996);
   U23997 : OAI22_X1 port map( A1 => n9107, A2 => n30591, B1 => n31054, B2 => 
                           n30585, ZN => n5997);
   U23998 : OAI22_X1 port map( A1 => n9102, A2 => n30591, B1 => n31057, B2 => 
                           n30585, ZN => n5998);
   U23999 : OAI22_X1 port map( A1 => n9097, A2 => n30591, B1 => n31060, B2 => 
                           n30585, ZN => n5999);
   U24000 : OAI22_X1 port map( A1 => n9092, A2 => n30591, B1 => n31063, B2 => 
                           n30585, ZN => n6000);
   U24001 : OAI22_X1 port map( A1 => n9087, A2 => n30591, B1 => n31066, B2 => 
                           n30585, ZN => n6001);
   U24002 : OAI22_X1 port map( A1 => n9082, A2 => n30591, B1 => n31069, B2 => 
                           n30585, ZN => n6002);
   U24003 : OAI22_X1 port map( A1 => n9077, A2 => n30591, B1 => n31072, B2 => 
                           n30585, ZN => n6003);
   U24004 : OAI22_X1 port map( A1 => n9072, A2 => n30591, B1 => n31075, B2 => 
                           n30585, ZN => n6004);
   U24005 : OAI22_X1 port map( A1 => n9067, A2 => n30591, B1 => n31078, B2 => 
                           n30585, ZN => n6005);
   U24006 : OAI22_X1 port map( A1 => n9062, A2 => n30591, B1 => n31081, B2 => 
                           n30585, ZN => n6006);
   U24007 : OAI22_X1 port map( A1 => n9057, A2 => n30591, B1 => n31084, B2 => 
                           n30585, ZN => n6007);
   U24008 : OAI22_X1 port map( A1 => n9052, A2 => n30592, B1 => n31087, B2 => 
                           n30585, ZN => n6008);
   U24009 : OAI22_X1 port map( A1 => n9047, A2 => n30592, B1 => n31090, B2 => 
                           n30586, ZN => n6009);
   U24010 : OAI22_X1 port map( A1 => n9042, A2 => n30592, B1 => n31093, B2 => 
                           n30586, ZN => n6010);
   U24011 : OAI22_X1 port map( A1 => n9037, A2 => n30592, B1 => n31096, B2 => 
                           n30586, ZN => n6011);
   U24012 : OAI22_X1 port map( A1 => n9032, A2 => n30592, B1 => n31099, B2 => 
                           n30586, ZN => n6012);
   U24013 : OAI22_X1 port map( A1 => n9027, A2 => n30592, B1 => n31102, B2 => 
                           n30586, ZN => n6013);
   U24014 : OAI22_X1 port map( A1 => n9022, A2 => n30592, B1 => n31105, B2 => 
                           n30586, ZN => n6014);
   U24015 : OAI22_X1 port map( A1 => n9017, A2 => n30592, B1 => n31108, B2 => 
                           n30586, ZN => n6015);
   U24016 : OAI22_X1 port map( A1 => n9012, A2 => n30592, B1 => n31111, B2 => 
                           n30586, ZN => n6016);
   U24017 : OAI22_X1 port map( A1 => n9007, A2 => n30592, B1 => n31114, B2 => 
                           n30586, ZN => n6017);
   U24018 : OAI22_X1 port map( A1 => n9002, A2 => n30592, B1 => n31117, B2 => 
                           n30586, ZN => n6018);
   U24019 : OAI22_X1 port map( A1 => n8997, A2 => n30592, B1 => n31120, B2 => 
                           n30586, ZN => n6019);
   U24020 : OAI22_X1 port map( A1 => n8992, A2 => n30593, B1 => n31123, B2 => 
                           n30586, ZN => n6020);
   U24021 : OAI22_X1 port map( A1 => n9995, A2 => n30604, B1 => n30982, B2 => 
                           n30595, ZN => n6037);
   U24022 : OAI22_X1 port map( A1 => n9990, A2 => n30604, B1 => n30985, B2 => 
                           n30595, ZN => n6038);
   U24023 : OAI22_X1 port map( A1 => n9985, A2 => n30604, B1 => n30988, B2 => 
                           n30595, ZN => n6039);
   U24024 : OAI22_X1 port map( A1 => n9980, A2 => n30604, B1 => n30991, B2 => 
                           n30595, ZN => n6040);
   U24025 : OAI22_X1 port map( A1 => n9975, A2 => n30604, B1 => n30994, B2 => 
                           n30595, ZN => n6041);
   U24026 : OAI22_X1 port map( A1 => n9970, A2 => n30603, B1 => n30997, B2 => 
                           n30595, ZN => n6042);
   U24027 : OAI22_X1 port map( A1 => n9965, A2 => n30603, B1 => n31000, B2 => 
                           n30595, ZN => n6043);
   U24028 : OAI22_X1 port map( A1 => n9960, A2 => n30603, B1 => n31003, B2 => 
                           n30595, ZN => n6044);
   U24029 : OAI22_X1 port map( A1 => n9955, A2 => n30603, B1 => n31006, B2 => 
                           n30595, ZN => n6045);
   U24030 : OAI22_X1 port map( A1 => n9950, A2 => n30603, B1 => n31009, B2 => 
                           n30595, ZN => n6046);
   U24031 : OAI22_X1 port map( A1 => n9945, A2 => n30603, B1 => n31012, B2 => 
                           n30595, ZN => n6047);
   U24032 : OAI22_X1 port map( A1 => n9940, A2 => n30603, B1 => n31015, B2 => 
                           n30595, ZN => n6048);
   U24033 : OAI22_X1 port map( A1 => n9935, A2 => n30603, B1 => n31018, B2 => 
                           n30596, ZN => n6049);
   U24034 : OAI22_X1 port map( A1 => n9930, A2 => n30603, B1 => n31021, B2 => 
                           n30596, ZN => n6050);
   U24035 : OAI22_X1 port map( A1 => n9925, A2 => n30603, B1 => n31024, B2 => 
                           n30596, ZN => n6051);
   U24036 : OAI22_X1 port map( A1 => n9920, A2 => n30603, B1 => n31027, B2 => 
                           n30596, ZN => n6052);
   U24037 : OAI22_X1 port map( A1 => n9915, A2 => n30603, B1 => n31030, B2 => 
                           n30596, ZN => n6053);
   U24038 : OAI22_X1 port map( A1 => n9910, A2 => n30602, B1 => n31033, B2 => 
                           n30596, ZN => n6054);
   U24039 : OAI22_X1 port map( A1 => n9905, A2 => n30602, B1 => n31036, B2 => 
                           n30596, ZN => n6055);
   U24040 : OAI22_X1 port map( A1 => n9900, A2 => n30602, B1 => n31039, B2 => 
                           n30596, ZN => n6056);
   U24041 : OAI22_X1 port map( A1 => n9895, A2 => n30602, B1 => n31042, B2 => 
                           n30596, ZN => n6057);
   U24042 : OAI22_X1 port map( A1 => n9890, A2 => n30602, B1 => n31045, B2 => 
                           n30596, ZN => n6058);
   U24043 : OAI22_X1 port map( A1 => n9885, A2 => n30602, B1 => n31048, B2 => 
                           n30596, ZN => n6059);
   U24044 : OAI22_X1 port map( A1 => n9880, A2 => n30602, B1 => n31051, B2 => 
                           n30596, ZN => n6060);
   U24045 : OAI22_X1 port map( A1 => n9875, A2 => n30602, B1 => n31054, B2 => 
                           n30597, ZN => n6061);
   U24046 : OAI22_X1 port map( A1 => n9870, A2 => n30602, B1 => n31057, B2 => 
                           n30597, ZN => n6062);
   U24047 : OAI22_X1 port map( A1 => n9865, A2 => n30602, B1 => n31060, B2 => 
                           n30597, ZN => n6063);
   U24048 : OAI22_X1 port map( A1 => n9860, A2 => n30602, B1 => n31063, B2 => 
                           n30597, ZN => n6064);
   U24049 : OAI22_X1 port map( A1 => n9855, A2 => n30601, B1 => n31066, B2 => 
                           n30597, ZN => n6065);
   U24050 : OAI22_X1 port map( A1 => n9850, A2 => n30601, B1 => n31069, B2 => 
                           n30597, ZN => n6066);
   U24051 : OAI22_X1 port map( A1 => n9845, A2 => n30601, B1 => n31072, B2 => 
                           n30597, ZN => n6067);
   U24052 : OAI22_X1 port map( A1 => n9840, A2 => n30601, B1 => n31075, B2 => 
                           n30597, ZN => n6068);
   U24053 : OAI22_X1 port map( A1 => n9835, A2 => n30601, B1 => n31078, B2 => 
                           n30597, ZN => n6069);
   U24054 : OAI22_X1 port map( A1 => n9830, A2 => n30601, B1 => n31081, B2 => 
                           n30597, ZN => n6070);
   U24055 : OAI22_X1 port map( A1 => n9825, A2 => n30601, B1 => n31084, B2 => 
                           n30597, ZN => n6071);
   U24056 : OAI22_X1 port map( A1 => n9820, A2 => n30601, B1 => n31087, B2 => 
                           n30597, ZN => n6072);
   U24057 : OAI22_X1 port map( A1 => n9815, A2 => n30601, B1 => n31090, B2 => 
                           n30598, ZN => n6073);
   U24058 : OAI22_X1 port map( A1 => n9810, A2 => n30601, B1 => n31093, B2 => 
                           n30598, ZN => n6074);
   U24059 : OAI22_X1 port map( A1 => n9805, A2 => n30601, B1 => n31096, B2 => 
                           n30598, ZN => n6075);
   U24060 : OAI22_X1 port map( A1 => n9800, A2 => n30601, B1 => n31099, B2 => 
                           n30598, ZN => n6076);
   U24061 : OAI22_X1 port map( A1 => n9795, A2 => n30600, B1 => n31102, B2 => 
                           n30598, ZN => n6077);
   U24062 : OAI22_X1 port map( A1 => n9790, A2 => n30600, B1 => n31105, B2 => 
                           n30598, ZN => n6078);
   U24063 : OAI22_X1 port map( A1 => n9785, A2 => n30600, B1 => n31108, B2 => 
                           n30598, ZN => n6079);
   U24064 : OAI22_X1 port map( A1 => n9780, A2 => n30600, B1 => n31111, B2 => 
                           n30598, ZN => n6080);
   U24065 : OAI22_X1 port map( A1 => n9775, A2 => n30600, B1 => n31114, B2 => 
                           n30598, ZN => n6081);
   U24066 : OAI22_X1 port map( A1 => n9770, A2 => n30600, B1 => n31117, B2 => 
                           n30598, ZN => n6082);
   U24067 : OAI22_X1 port map( A1 => n9765, A2 => n30600, B1 => n31120, B2 => 
                           n30598, ZN => n6083);
   U24068 : OAI22_X1 port map( A1 => n9760, A2 => n30600, B1 => n31123, B2 => 
                           n30598, ZN => n6084);
   U24069 : OAI22_X1 port map( A1 => n30614, A2 => n26233, B1 => n30946, B2 => 
                           n30606, ZN => n6089);
   U24070 : OAI22_X1 port map( A1 => n30614, A2 => n26232, B1 => n30949, B2 => 
                           n30606, ZN => n6090);
   U24071 : OAI22_X1 port map( A1 => n30614, A2 => n26231, B1 => n30952, B2 => 
                           n30606, ZN => n6091);
   U24072 : OAI22_X1 port map( A1 => n30614, A2 => n26230, B1 => n30955, B2 => 
                           n30606, ZN => n6092);
   U24073 : OAI22_X1 port map( A1 => n30614, A2 => n26229, B1 => n30958, B2 => 
                           n30606, ZN => n6093);
   U24074 : OAI22_X1 port map( A1 => n30614, A2 => n26228, B1 => n30961, B2 => 
                           n30606, ZN => n6094);
   U24075 : OAI22_X1 port map( A1 => n30614, A2 => n26227, B1 => n30964, B2 => 
                           n30606, ZN => n6095);
   U24076 : OAI22_X1 port map( A1 => n30614, A2 => n26226, B1 => n30967, B2 => 
                           n30606, ZN => n6096);
   U24077 : OAI22_X1 port map( A1 => n30614, A2 => n26225, B1 => n30970, B2 => 
                           n30606, ZN => n6097);
   U24078 : OAI22_X1 port map( A1 => n30614, A2 => n26224, B1 => n30973, B2 => 
                           n30606, ZN => n6098);
   U24079 : OAI22_X1 port map( A1 => n30614, A2 => n26223, B1 => n30976, B2 => 
                           n30606, ZN => n6099);
   U24080 : OAI22_X1 port map( A1 => n30614, A2 => n26222, B1 => n30979, B2 => 
                           n30606, ZN => n6100);
   U24081 : OAI22_X1 port map( A1 => n30615, A2 => n26221, B1 => n30982, B2 => 
                           n30607, ZN => n6101);
   U24082 : OAI22_X1 port map( A1 => n30615, A2 => n26220, B1 => n30985, B2 => 
                           n30607, ZN => n6102);
   U24083 : OAI22_X1 port map( A1 => n30615, A2 => n26219, B1 => n30988, B2 => 
                           n30607, ZN => n6103);
   U24084 : OAI22_X1 port map( A1 => n30615, A2 => n26218, B1 => n30991, B2 => 
                           n30607, ZN => n6104);
   U24085 : OAI22_X1 port map( A1 => n30615, A2 => n26217, B1 => n30994, B2 => 
                           n30607, ZN => n6105);
   U24086 : OAI22_X1 port map( A1 => n30615, A2 => n26216, B1 => n30997, B2 => 
                           n30607, ZN => n6106);
   U24087 : OAI22_X1 port map( A1 => n30615, A2 => n26215, B1 => n31000, B2 => 
                           n30607, ZN => n6107);
   U24088 : OAI22_X1 port map( A1 => n30615, A2 => n26214, B1 => n31003, B2 => 
                           n30607, ZN => n6108);
   U24089 : OAI22_X1 port map( A1 => n30615, A2 => n26213, B1 => n31006, B2 => 
                           n30607, ZN => n6109);
   U24090 : OAI22_X1 port map( A1 => n30615, A2 => n26212, B1 => n31009, B2 => 
                           n30607, ZN => n6110);
   U24091 : OAI22_X1 port map( A1 => n30615, A2 => n26211, B1 => n31012, B2 => 
                           n30607, ZN => n6111);
   U24092 : OAI22_X1 port map( A1 => n30615, A2 => n26210, B1 => n31015, B2 => 
                           n30607, ZN => n6112);
   U24093 : OAI22_X1 port map( A1 => n30615, A2 => n26209, B1 => n31018, B2 => 
                           n30608, ZN => n6113);
   U24094 : OAI22_X1 port map( A1 => n30616, A2 => n26208, B1 => n31021, B2 => 
                           n30608, ZN => n6114);
   U24095 : OAI22_X1 port map( A1 => n30616, A2 => n26207, B1 => n31024, B2 => 
                           n30608, ZN => n6115);
   U24096 : OAI22_X1 port map( A1 => n30616, A2 => n26206, B1 => n31027, B2 => 
                           n30608, ZN => n6116);
   U24097 : OAI22_X1 port map( A1 => n30616, A2 => n26205, B1 => n31030, B2 => 
                           n30608, ZN => n6117);
   U24098 : OAI22_X1 port map( A1 => n30616, A2 => n26204, B1 => n31033, B2 => 
                           n30608, ZN => n6118);
   U24099 : OAI22_X1 port map( A1 => n30616, A2 => n26203, B1 => n31036, B2 => 
                           n30608, ZN => n6119);
   U24100 : OAI22_X1 port map( A1 => n30616, A2 => n26202, B1 => n31039, B2 => 
                           n30608, ZN => n6120);
   U24101 : OAI22_X1 port map( A1 => n30616, A2 => n26201, B1 => n31042, B2 => 
                           n30608, ZN => n6121);
   U24102 : OAI22_X1 port map( A1 => n30616, A2 => n26200, B1 => n31045, B2 => 
                           n30608, ZN => n6122);
   U24103 : OAI22_X1 port map( A1 => n30616, A2 => n26199, B1 => n31048, B2 => 
                           n30608, ZN => n6123);
   U24104 : OAI22_X1 port map( A1 => n30616, A2 => n26198, B1 => n31051, B2 => 
                           n30608, ZN => n6124);
   U24105 : OAI22_X1 port map( A1 => n30616, A2 => n26197, B1 => n31054, B2 => 
                           n30609, ZN => n6125);
   U24106 : OAI22_X1 port map( A1 => n30616, A2 => n26196, B1 => n31057, B2 => 
                           n30609, ZN => n6126);
   U24107 : OAI22_X1 port map( A1 => n30617, A2 => n26195, B1 => n31060, B2 => 
                           n30609, ZN => n6127);
   U24108 : OAI22_X1 port map( A1 => n30617, A2 => n26194, B1 => n31063, B2 => 
                           n30609, ZN => n6128);
   U24109 : OAI22_X1 port map( A1 => n30617, A2 => n26193, B1 => n31066, B2 => 
                           n30609, ZN => n6129);
   U24110 : OAI22_X1 port map( A1 => n30617, A2 => n26192, B1 => n31069, B2 => 
                           n30609, ZN => n6130);
   U24111 : OAI22_X1 port map( A1 => n30617, A2 => n26191, B1 => n31072, B2 => 
                           n30609, ZN => n6131);
   U24112 : OAI22_X1 port map( A1 => n30617, A2 => n26190, B1 => n31075, B2 => 
                           n30609, ZN => n6132);
   U24113 : OAI22_X1 port map( A1 => n30617, A2 => n26189, B1 => n31078, B2 => 
                           n30609, ZN => n6133);
   U24114 : OAI22_X1 port map( A1 => n30617, A2 => n26188, B1 => n31081, B2 => 
                           n30609, ZN => n6134);
   U24115 : OAI22_X1 port map( A1 => n30617, A2 => n26187, B1 => n31084, B2 => 
                           n30609, ZN => n6135);
   U24116 : OAI22_X1 port map( A1 => n30617, A2 => n26186, B1 => n31087, B2 => 
                           n30609, ZN => n6136);
   U24117 : OAI22_X1 port map( A1 => n30617, A2 => n26185, B1 => n31090, B2 => 
                           n30610, ZN => n6137);
   U24118 : OAI22_X1 port map( A1 => n30617, A2 => n26184, B1 => n31093, B2 => 
                           n30610, ZN => n6138);
   U24119 : OAI22_X1 port map( A1 => n30617, A2 => n26183, B1 => n31096, B2 => 
                           n30610, ZN => n6139);
   U24120 : OAI22_X1 port map( A1 => n30618, A2 => n26182, B1 => n31099, B2 => 
                           n30610, ZN => n6140);
   U24121 : OAI22_X1 port map( A1 => n30618, A2 => n26181, B1 => n31102, B2 => 
                           n30610, ZN => n6141);
   U24122 : OAI22_X1 port map( A1 => n30618, A2 => n26180, B1 => n31105, B2 => 
                           n30610, ZN => n6142);
   U24123 : OAI22_X1 port map( A1 => n30618, A2 => n26179, B1 => n31108, B2 => 
                           n30610, ZN => n6143);
   U24124 : OAI22_X1 port map( A1 => n30618, A2 => n26178, B1 => n31111, B2 => 
                           n30610, ZN => n6144);
   U24125 : OAI22_X1 port map( A1 => n30618, A2 => n26177, B1 => n31114, B2 => 
                           n30610, ZN => n6145);
   U24126 : OAI22_X1 port map( A1 => n30618, A2 => n26176, B1 => n31117, B2 => 
                           n30610, ZN => n6146);
   U24127 : OAI22_X1 port map( A1 => n30618, A2 => n26175, B1 => n31120, B2 => 
                           n30610, ZN => n6147);
   U24128 : OAI22_X1 port map( A1 => n30618, A2 => n26174, B1 => n31123, B2 => 
                           n30610, ZN => n6148);
   U24129 : OAI22_X1 port map( A1 => n30851, A2 => n25586, B1 => n30945, B2 => 
                           n30843, ZN => n7305);
   U24130 : OAI22_X1 port map( A1 => n30851, A2 => n25585, B1 => n30948, B2 => 
                           n30843, ZN => n7306);
   U24131 : OAI22_X1 port map( A1 => n30851, A2 => n25584, B1 => n30951, B2 => 
                           n30843, ZN => n7307);
   U24132 : OAI22_X1 port map( A1 => n30851, A2 => n25583, B1 => n30954, B2 => 
                           n30843, ZN => n7308);
   U24133 : OAI22_X1 port map( A1 => n30851, A2 => n25582, B1 => n30957, B2 => 
                           n30843, ZN => n7309);
   U24134 : OAI22_X1 port map( A1 => n30851, A2 => n25581, B1 => n30960, B2 => 
                           n30843, ZN => n7310);
   U24135 : OAI22_X1 port map( A1 => n30851, A2 => n25580, B1 => n30963, B2 => 
                           n30843, ZN => n7311);
   U24136 : OAI22_X1 port map( A1 => n30851, A2 => n25579, B1 => n30966, B2 => 
                           n30843, ZN => n7312);
   U24137 : OAI22_X1 port map( A1 => n30851, A2 => n25578, B1 => n30969, B2 => 
                           n30843, ZN => n7313);
   U24138 : OAI22_X1 port map( A1 => n30851, A2 => n25577, B1 => n30972, B2 => 
                           n30843, ZN => n7314);
   U24139 : OAI22_X1 port map( A1 => n30851, A2 => n25576, B1 => n30975, B2 => 
                           n30843, ZN => n7315);
   U24140 : OAI22_X1 port map( A1 => n30851, A2 => n25575, B1 => n30978, B2 => 
                           n30843, ZN => n7316);
   U24141 : OAI22_X1 port map( A1 => n30852, A2 => n25574, B1 => n30981, B2 => 
                           n30844, ZN => n7317);
   U24142 : OAI22_X1 port map( A1 => n30852, A2 => n25573, B1 => n30984, B2 => 
                           n30844, ZN => n7318);
   U24143 : OAI22_X1 port map( A1 => n30852, A2 => n25572, B1 => n30987, B2 => 
                           n30844, ZN => n7319);
   U24144 : OAI22_X1 port map( A1 => n30852, A2 => n25571, B1 => n30990, B2 => 
                           n30844, ZN => n7320);
   U24145 : OAI22_X1 port map( A1 => n30852, A2 => n25570, B1 => n30993, B2 => 
                           n30844, ZN => n7321);
   U24146 : OAI22_X1 port map( A1 => n30852, A2 => n25569, B1 => n30996, B2 => 
                           n30844, ZN => n7322);
   U24147 : OAI22_X1 port map( A1 => n30852, A2 => n25568, B1 => n30999, B2 => 
                           n30844, ZN => n7323);
   U24148 : OAI22_X1 port map( A1 => n30852, A2 => n25567, B1 => n31002, B2 => 
                           n30844, ZN => n7324);
   U24149 : OAI22_X1 port map( A1 => n30852, A2 => n25566, B1 => n31005, B2 => 
                           n30844, ZN => n7325);
   U24150 : OAI22_X1 port map( A1 => n30852, A2 => n25565, B1 => n31008, B2 => 
                           n30844, ZN => n7326);
   U24151 : OAI22_X1 port map( A1 => n30852, A2 => n25564, B1 => n31011, B2 => 
                           n30844, ZN => n7327);
   U24152 : OAI22_X1 port map( A1 => n30852, A2 => n25563, B1 => n31014, B2 => 
                           n30844, ZN => n7328);
   U24153 : OAI22_X1 port map( A1 => n30852, A2 => n25562, B1 => n31017, B2 => 
                           n30845, ZN => n7329);
   U24154 : OAI22_X1 port map( A1 => n30853, A2 => n25561, B1 => n31020, B2 => 
                           n30845, ZN => n7330);
   U24155 : OAI22_X1 port map( A1 => n30853, A2 => n25560, B1 => n31023, B2 => 
                           n30845, ZN => n7331);
   U24156 : OAI22_X1 port map( A1 => n30853, A2 => n25559, B1 => n31026, B2 => 
                           n30845, ZN => n7332);
   U24157 : OAI22_X1 port map( A1 => n30853, A2 => n25558, B1 => n31029, B2 => 
                           n30845, ZN => n7333);
   U24158 : OAI22_X1 port map( A1 => n30853, A2 => n25557, B1 => n31032, B2 => 
                           n30845, ZN => n7334);
   U24159 : OAI22_X1 port map( A1 => n30853, A2 => n25556, B1 => n31035, B2 => 
                           n30845, ZN => n7335);
   U24160 : OAI22_X1 port map( A1 => n30853, A2 => n25555, B1 => n31038, B2 => 
                           n30845, ZN => n7336);
   U24161 : OAI22_X1 port map( A1 => n30853, A2 => n25554, B1 => n31041, B2 => 
                           n30845, ZN => n7337);
   U24162 : OAI22_X1 port map( A1 => n30853, A2 => n25553, B1 => n31044, B2 => 
                           n30845, ZN => n7338);
   U24163 : OAI22_X1 port map( A1 => n30853, A2 => n25552, B1 => n31047, B2 => 
                           n30845, ZN => n7339);
   U24164 : OAI22_X1 port map( A1 => n30853, A2 => n25551, B1 => n31050, B2 => 
                           n30845, ZN => n7340);
   U24165 : OAI22_X1 port map( A1 => n30853, A2 => n25550, B1 => n31053, B2 => 
                           n30846, ZN => n7341);
   U24166 : OAI22_X1 port map( A1 => n30853, A2 => n25549, B1 => n31056, B2 => 
                           n30846, ZN => n7342);
   U24167 : OAI22_X1 port map( A1 => n30854, A2 => n25548, B1 => n31059, B2 => 
                           n30846, ZN => n7343);
   U24168 : OAI22_X1 port map( A1 => n30854, A2 => n25547, B1 => n31062, B2 => 
                           n30846, ZN => n7344);
   U24169 : OAI22_X1 port map( A1 => n30854, A2 => n25546, B1 => n31065, B2 => 
                           n30846, ZN => n7345);
   U24170 : OAI22_X1 port map( A1 => n30854, A2 => n25545, B1 => n31068, B2 => 
                           n30846, ZN => n7346);
   U24171 : OAI22_X1 port map( A1 => n30854, A2 => n25544, B1 => n31071, B2 => 
                           n30846, ZN => n7347);
   U24172 : OAI22_X1 port map( A1 => n30854, A2 => n25543, B1 => n31074, B2 => 
                           n30846, ZN => n7348);
   U24173 : OAI22_X1 port map( A1 => n30854, A2 => n25542, B1 => n31077, B2 => 
                           n30846, ZN => n7349);
   U24174 : OAI22_X1 port map( A1 => n30854, A2 => n25541, B1 => n31080, B2 => 
                           n30846, ZN => n7350);
   U24175 : OAI22_X1 port map( A1 => n30854, A2 => n25540, B1 => n31083, B2 => 
                           n30846, ZN => n7351);
   U24176 : OAI22_X1 port map( A1 => n30854, A2 => n25539, B1 => n31086, B2 => 
                           n30846, ZN => n7352);
   U24177 : OAI22_X1 port map( A1 => n30854, A2 => n25538, B1 => n31089, B2 => 
                           n30847, ZN => n7353);
   U24178 : OAI22_X1 port map( A1 => n30854, A2 => n25537, B1 => n31092, B2 => 
                           n30847, ZN => n7354);
   U24179 : OAI22_X1 port map( A1 => n30854, A2 => n25536, B1 => n31095, B2 => 
                           n30847, ZN => n7355);
   U24180 : OAI22_X1 port map( A1 => n30855, A2 => n25535, B1 => n31098, B2 => 
                           n30847, ZN => n7356);
   U24181 : OAI22_X1 port map( A1 => n30855, A2 => n25534, B1 => n31101, B2 => 
                           n30847, ZN => n7357);
   U24182 : OAI22_X1 port map( A1 => n30855, A2 => n25533, B1 => n31104, B2 => 
                           n30847, ZN => n7358);
   U24183 : OAI22_X1 port map( A1 => n30855, A2 => n25532, B1 => n31107, B2 => 
                           n30847, ZN => n7359);
   U24184 : OAI22_X1 port map( A1 => n30855, A2 => n25531, B1 => n31110, B2 => 
                           n30847, ZN => n7360);
   U24185 : OAI22_X1 port map( A1 => n30855, A2 => n25530, B1 => n31113, B2 => 
                           n30847, ZN => n7361);
   U24186 : OAI22_X1 port map( A1 => n30855, A2 => n25529, B1 => n31116, B2 => 
                           n30847, ZN => n7362);
   U24187 : OAI22_X1 port map( A1 => n30855, A2 => n25528, B1 => n31119, B2 => 
                           n30847, ZN => n7363);
   U24188 : OAI22_X1 port map( A1 => n30855, A2 => n25527, B1 => n31122, B2 => 
                           n30847, ZN => n7364);
   U24189 : OAI22_X1 port map( A1 => n17836, A2 => n30774, B1 => n30945, B2 => 
                           n30768, ZN => n6921);
   U24190 : OAI22_X1 port map( A1 => n17835, A2 => n30774, B1 => n30948, B2 => 
                           n30768, ZN => n6922);
   U24191 : OAI22_X1 port map( A1 => n17834, A2 => n30774, B1 => n30951, B2 => 
                           n30768, ZN => n6923);
   U24192 : OAI22_X1 port map( A1 => n17833, A2 => n30774, B1 => n30954, B2 => 
                           n30768, ZN => n6924);
   U24193 : OAI22_X1 port map( A1 => n17832, A2 => n30774, B1 => n30957, B2 => 
                           n30768, ZN => n6925);
   U24194 : OAI22_X1 port map( A1 => n17831, A2 => n30774, B1 => n30960, B2 => 
                           n30768, ZN => n6926);
   U24195 : OAI22_X1 port map( A1 => n17830, A2 => n30774, B1 => n30963, B2 => 
                           n30768, ZN => n6927);
   U24196 : OAI22_X1 port map( A1 => n17829, A2 => n30774, B1 => n30966, B2 => 
                           n30768, ZN => n6928);
   U24197 : OAI22_X1 port map( A1 => n17828, A2 => n30774, B1 => n30969, B2 => 
                           n30768, ZN => n6929);
   U24198 : OAI22_X1 port map( A1 => n17827, A2 => n30774, B1 => n30972, B2 => 
                           n30768, ZN => n6930);
   U24199 : OAI22_X1 port map( A1 => n17826, A2 => n30774, B1 => n30975, B2 => 
                           n30768, ZN => n6931);
   U24200 : OAI22_X1 port map( A1 => n17825, A2 => n30775, B1 => n30978, B2 => 
                           n30768, ZN => n6932);
   U24201 : OAI22_X1 port map( A1 => n17824, A2 => n30775, B1 => n30981, B2 => 
                           n30769, ZN => n6933);
   U24202 : OAI22_X1 port map( A1 => n17823, A2 => n30775, B1 => n30984, B2 => 
                           n30769, ZN => n6934);
   U24203 : OAI22_X1 port map( A1 => n17822, A2 => n30775, B1 => n30987, B2 => 
                           n30769, ZN => n6935);
   U24204 : OAI22_X1 port map( A1 => n17821, A2 => n30775, B1 => n30990, B2 => 
                           n30769, ZN => n6936);
   U24205 : OAI22_X1 port map( A1 => n17820, A2 => n30775, B1 => n30993, B2 => 
                           n30769, ZN => n6937);
   U24206 : OAI22_X1 port map( A1 => n17819, A2 => n30775, B1 => n30996, B2 => 
                           n30769, ZN => n6938);
   U24207 : OAI22_X1 port map( A1 => n17818, A2 => n30775, B1 => n30999, B2 => 
                           n30769, ZN => n6939);
   U24208 : OAI22_X1 port map( A1 => n17817, A2 => n30775, B1 => n31002, B2 => 
                           n30769, ZN => n6940);
   U24209 : OAI22_X1 port map( A1 => n17816, A2 => n30775, B1 => n31005, B2 => 
                           n30769, ZN => n6941);
   U24210 : OAI22_X1 port map( A1 => n17815, A2 => n30775, B1 => n31008, B2 => 
                           n30769, ZN => n6942);
   U24211 : OAI22_X1 port map( A1 => n17814, A2 => n30775, B1 => n31011, B2 => 
                           n30769, ZN => n6943);
   U24212 : OAI22_X1 port map( A1 => n17813, A2 => n30776, B1 => n31014, B2 => 
                           n30769, ZN => n6944);
   U24213 : OAI22_X1 port map( A1 => n17812, A2 => n30776, B1 => n31017, B2 => 
                           n30770, ZN => n6945);
   U24214 : OAI22_X1 port map( A1 => n17811, A2 => n30776, B1 => n31020, B2 => 
                           n30770, ZN => n6946);
   U24215 : OAI22_X1 port map( A1 => n17810, A2 => n30776, B1 => n31023, B2 => 
                           n30770, ZN => n6947);
   U24216 : OAI22_X1 port map( A1 => n17809, A2 => n30776, B1 => n31026, B2 => 
                           n30770, ZN => n6948);
   U24217 : OAI22_X1 port map( A1 => n17808, A2 => n30776, B1 => n31029, B2 => 
                           n30770, ZN => n6949);
   U24218 : OAI22_X1 port map( A1 => n17807, A2 => n30776, B1 => n31032, B2 => 
                           n30770, ZN => n6950);
   U24219 : OAI22_X1 port map( A1 => n17806, A2 => n30776, B1 => n31035, B2 => 
                           n30770, ZN => n6951);
   U24220 : OAI22_X1 port map( A1 => n17805, A2 => n30776, B1 => n31038, B2 => 
                           n30770, ZN => n6952);
   U24221 : OAI22_X1 port map( A1 => n17804, A2 => n30776, B1 => n31041, B2 => 
                           n30770, ZN => n6953);
   U24222 : OAI22_X1 port map( A1 => n17803, A2 => n30776, B1 => n31044, B2 => 
                           n30770, ZN => n6954);
   U24223 : OAI22_X1 port map( A1 => n17802, A2 => n30776, B1 => n31047, B2 => 
                           n30770, ZN => n6955);
   U24224 : OAI22_X1 port map( A1 => n17801, A2 => n30777, B1 => n31050, B2 => 
                           n30770, ZN => n6956);
   U24225 : OAI22_X1 port map( A1 => n17800, A2 => n30777, B1 => n31053, B2 => 
                           n30771, ZN => n6957);
   U24226 : OAI22_X1 port map( A1 => n17799, A2 => n30777, B1 => n31056, B2 => 
                           n30771, ZN => n6958);
   U24227 : OAI22_X1 port map( A1 => n17798, A2 => n30777, B1 => n31059, B2 => 
                           n30771, ZN => n6959);
   U24228 : OAI22_X1 port map( A1 => n17797, A2 => n30777, B1 => n31062, B2 => 
                           n30771, ZN => n6960);
   U24229 : OAI22_X1 port map( A1 => n17796, A2 => n30777, B1 => n31065, B2 => 
                           n30771, ZN => n6961);
   U24230 : OAI22_X1 port map( A1 => n17795, A2 => n30777, B1 => n31068, B2 => 
                           n30771, ZN => n6962);
   U24231 : OAI22_X1 port map( A1 => n17794, A2 => n30777, B1 => n31071, B2 => 
                           n30771, ZN => n6963);
   U24232 : OAI22_X1 port map( A1 => n17793, A2 => n30777, B1 => n31074, B2 => 
                           n30771, ZN => n6964);
   U24233 : OAI22_X1 port map( A1 => n17792, A2 => n30777, B1 => n31077, B2 => 
                           n30771, ZN => n6965);
   U24234 : OAI22_X1 port map( A1 => n17791, A2 => n30777, B1 => n31080, B2 => 
                           n30771, ZN => n6966);
   U24235 : OAI22_X1 port map( A1 => n17790, A2 => n30777, B1 => n31083, B2 => 
                           n30771, ZN => n6967);
   U24236 : OAI22_X1 port map( A1 => n17789, A2 => n30778, B1 => n31086, B2 => 
                           n30771, ZN => n6968);
   U24237 : OAI22_X1 port map( A1 => n17788, A2 => n30778, B1 => n31089, B2 => 
                           n30772, ZN => n6969);
   U24238 : OAI22_X1 port map( A1 => n17787, A2 => n30778, B1 => n31092, B2 => 
                           n30772, ZN => n6970);
   U24239 : OAI22_X1 port map( A1 => n17786, A2 => n30778, B1 => n31095, B2 => 
                           n30772, ZN => n6971);
   U24240 : OAI22_X1 port map( A1 => n17785, A2 => n30778, B1 => n31098, B2 => 
                           n30772, ZN => n6972);
   U24241 : OAI22_X1 port map( A1 => n17784, A2 => n30778, B1 => n31101, B2 => 
                           n30772, ZN => n6973);
   U24242 : OAI22_X1 port map( A1 => n17783, A2 => n30778, B1 => n31104, B2 => 
                           n30772, ZN => n6974);
   U24243 : OAI22_X1 port map( A1 => n17782, A2 => n30778, B1 => n31107, B2 => 
                           n30772, ZN => n6975);
   U24244 : OAI22_X1 port map( A1 => n17781, A2 => n30778, B1 => n31110, B2 => 
                           n30772, ZN => n6976);
   U24245 : OAI22_X1 port map( A1 => n17780, A2 => n30778, B1 => n31113, B2 => 
                           n30772, ZN => n6977);
   U24246 : OAI22_X1 port map( A1 => n17779, A2 => n30778, B1 => n31116, B2 => 
                           n30772, ZN => n6978);
   U24247 : OAI22_X1 port map( A1 => n17778, A2 => n30778, B1 => n31119, B2 => 
                           n30772, ZN => n6979);
   U24248 : OAI22_X1 port map( A1 => n17777, A2 => n30779, B1 => n31122, B2 => 
                           n30772, ZN => n6980);
   U24249 : OAI22_X1 port map( A1 => n30927, A2 => n25301, B1 => n30944, B2 => 
                           n30919, ZN => n7689);
   U24250 : OAI22_X1 port map( A1 => n30927, A2 => n25300, B1 => n30947, B2 => 
                           n30919, ZN => n7690);
   U24251 : OAI22_X1 port map( A1 => n30927, A2 => n25299, B1 => n30950, B2 => 
                           n30919, ZN => n7691);
   U24252 : OAI22_X1 port map( A1 => n30927, A2 => n25298, B1 => n30953, B2 => 
                           n30919, ZN => n7692);
   U24253 : OAI22_X1 port map( A1 => n30927, A2 => n25297, B1 => n30956, B2 => 
                           n30919, ZN => n7693);
   U24254 : OAI22_X1 port map( A1 => n30927, A2 => n25296, B1 => n30959, B2 => 
                           n30919, ZN => n7694);
   U24255 : OAI22_X1 port map( A1 => n30927, A2 => n25295, B1 => n30962, B2 => 
                           n30919, ZN => n7695);
   U24256 : OAI22_X1 port map( A1 => n30927, A2 => n25294, B1 => n30965, B2 => 
                           n30919, ZN => n7696);
   U24257 : OAI22_X1 port map( A1 => n30927, A2 => n25293, B1 => n30968, B2 => 
                           n30919, ZN => n7697);
   U24258 : OAI22_X1 port map( A1 => n30927, A2 => n25292, B1 => n30971, B2 => 
                           n30919, ZN => n7698);
   U24259 : OAI22_X1 port map( A1 => n30927, A2 => n25291, B1 => n30974, B2 => 
                           n30919, ZN => n7699);
   U24260 : OAI22_X1 port map( A1 => n30927, A2 => n25290, B1 => n30977, B2 => 
                           n30919, ZN => n7700);
   U24261 : OAI22_X1 port map( A1 => n30928, A2 => n25289, B1 => n30980, B2 => 
                           n30920, ZN => n7701);
   U24262 : OAI22_X1 port map( A1 => n30928, A2 => n25288, B1 => n30983, B2 => 
                           n30920, ZN => n7702);
   U24263 : OAI22_X1 port map( A1 => n30928, A2 => n25287, B1 => n30986, B2 => 
                           n30920, ZN => n7703);
   U24264 : OAI22_X1 port map( A1 => n30928, A2 => n25286, B1 => n30989, B2 => 
                           n30920, ZN => n7704);
   U24265 : OAI22_X1 port map( A1 => n30928, A2 => n25285, B1 => n30992, B2 => 
                           n30920, ZN => n7705);
   U24266 : OAI22_X1 port map( A1 => n30928, A2 => n25284, B1 => n30995, B2 => 
                           n30920, ZN => n7706);
   U24267 : OAI22_X1 port map( A1 => n30928, A2 => n25283, B1 => n30998, B2 => 
                           n30920, ZN => n7707);
   U24268 : OAI22_X1 port map( A1 => n30928, A2 => n25282, B1 => n31001, B2 => 
                           n30920, ZN => n7708);
   U24269 : OAI22_X1 port map( A1 => n30928, A2 => n25281, B1 => n31004, B2 => 
                           n30920, ZN => n7709);
   U24270 : OAI22_X1 port map( A1 => n30928, A2 => n25280, B1 => n31007, B2 => 
                           n30920, ZN => n7710);
   U24271 : OAI22_X1 port map( A1 => n30928, A2 => n25279, B1 => n31010, B2 => 
                           n30920, ZN => n7711);
   U24272 : OAI22_X1 port map( A1 => n30928, A2 => n25278, B1 => n31013, B2 => 
                           n30920, ZN => n7712);
   U24273 : OAI22_X1 port map( A1 => n30928, A2 => n25277, B1 => n31016, B2 => 
                           n30921, ZN => n7713);
   U24274 : OAI22_X1 port map( A1 => n30929, A2 => n25276, B1 => n31019, B2 => 
                           n30921, ZN => n7714);
   U24275 : OAI22_X1 port map( A1 => n30929, A2 => n25275, B1 => n31022, B2 => 
                           n30921, ZN => n7715);
   U24276 : OAI22_X1 port map( A1 => n30929, A2 => n25274, B1 => n31025, B2 => 
                           n30921, ZN => n7716);
   U24277 : OAI22_X1 port map( A1 => n30929, A2 => n25273, B1 => n31028, B2 => 
                           n30921, ZN => n7717);
   U24278 : OAI22_X1 port map( A1 => n30929, A2 => n25272, B1 => n31031, B2 => 
                           n30921, ZN => n7718);
   U24279 : OAI22_X1 port map( A1 => n30929, A2 => n25271, B1 => n31034, B2 => 
                           n30921, ZN => n7719);
   U24280 : OAI22_X1 port map( A1 => n30929, A2 => n25270, B1 => n31037, B2 => 
                           n30921, ZN => n7720);
   U24281 : OAI22_X1 port map( A1 => n30929, A2 => n25269, B1 => n31040, B2 => 
                           n30921, ZN => n7721);
   U24282 : OAI22_X1 port map( A1 => n30929, A2 => n25268, B1 => n31043, B2 => 
                           n30921, ZN => n7722);
   U24283 : OAI22_X1 port map( A1 => n30929, A2 => n25267, B1 => n31046, B2 => 
                           n30921, ZN => n7723);
   U24284 : OAI22_X1 port map( A1 => n30929, A2 => n25266, B1 => n31049, B2 => 
                           n30921, ZN => n7724);
   U24285 : OAI22_X1 port map( A1 => n30929, A2 => n25265, B1 => n31052, B2 => 
                           n30922, ZN => n7725);
   U24286 : OAI22_X1 port map( A1 => n30929, A2 => n25264, B1 => n31055, B2 => 
                           n30922, ZN => n7726);
   U24287 : OAI22_X1 port map( A1 => n30930, A2 => n25263, B1 => n31058, B2 => 
                           n30922, ZN => n7727);
   U24288 : OAI22_X1 port map( A1 => n30930, A2 => n25262, B1 => n31061, B2 => 
                           n30922, ZN => n7728);
   U24289 : OAI22_X1 port map( A1 => n30930, A2 => n25261, B1 => n31064, B2 => 
                           n30922, ZN => n7729);
   U24290 : OAI22_X1 port map( A1 => n30930, A2 => n25260, B1 => n31067, B2 => 
                           n30922, ZN => n7730);
   U24291 : OAI22_X1 port map( A1 => n30930, A2 => n25259, B1 => n31070, B2 => 
                           n30922, ZN => n7731);
   U24292 : OAI22_X1 port map( A1 => n30930, A2 => n25258, B1 => n31073, B2 => 
                           n30922, ZN => n7732);
   U24293 : OAI22_X1 port map( A1 => n30930, A2 => n25257, B1 => n31076, B2 => 
                           n30922, ZN => n7733);
   U24294 : OAI22_X1 port map( A1 => n30930, A2 => n25256, B1 => n31079, B2 => 
                           n30922, ZN => n7734);
   U24295 : OAI22_X1 port map( A1 => n30930, A2 => n25255, B1 => n31082, B2 => 
                           n30922, ZN => n7735);
   U24296 : OAI22_X1 port map( A1 => n30930, A2 => n25254, B1 => n31085, B2 => 
                           n30922, ZN => n7736);
   U24297 : OAI22_X1 port map( A1 => n30930, A2 => n25253, B1 => n31088, B2 => 
                           n30923, ZN => n7737);
   U24298 : OAI22_X1 port map( A1 => n30930, A2 => n25252, B1 => n31091, B2 => 
                           n30923, ZN => n7738);
   U24299 : OAI22_X1 port map( A1 => n30930, A2 => n25251, B1 => n31094, B2 => 
                           n30923, ZN => n7739);
   U24300 : OAI22_X1 port map( A1 => n30931, A2 => n25250, B1 => n31097, B2 => 
                           n30923, ZN => n7740);
   U24301 : OAI22_X1 port map( A1 => n30931, A2 => n25249, B1 => n31100, B2 => 
                           n30923, ZN => n7741);
   U24302 : OAI22_X1 port map( A1 => n30931, A2 => n25248, B1 => n31103, B2 => 
                           n30923, ZN => n7742);
   U24303 : OAI22_X1 port map( A1 => n30931, A2 => n25247, B1 => n31106, B2 => 
                           n30923, ZN => n7743);
   U24304 : OAI22_X1 port map( A1 => n30931, A2 => n25246, B1 => n31109, B2 => 
                           n30923, ZN => n7744);
   U24305 : OAI22_X1 port map( A1 => n30931, A2 => n25245, B1 => n31112, B2 => 
                           n30923, ZN => n7745);
   U24306 : OAI22_X1 port map( A1 => n30931, A2 => n25244, B1 => n31115, B2 => 
                           n30923, ZN => n7746);
   U24307 : OAI22_X1 port map( A1 => n30931, A2 => n25243, B1 => n31118, B2 => 
                           n30923, ZN => n7747);
   U24308 : OAI22_X1 port map( A1 => n30931, A2 => n25242, B1 => n31121, B2 => 
                           n30923, ZN => n7748);
   U24309 : OAI22_X1 port map( A1 => n30877, A2 => n25450, B1 => n30944, B2 => 
                           n30869, ZN => n7433);
   U24310 : OAI22_X1 port map( A1 => n30877, A2 => n25449, B1 => n30947, B2 => 
                           n30869, ZN => n7434);
   U24311 : OAI22_X1 port map( A1 => n30877, A2 => n25448, B1 => n30950, B2 => 
                           n30869, ZN => n7435);
   U24312 : OAI22_X1 port map( A1 => n30877, A2 => n25447, B1 => n30953, B2 => 
                           n30869, ZN => n7436);
   U24313 : OAI22_X1 port map( A1 => n30877, A2 => n25446, B1 => n30956, B2 => 
                           n30869, ZN => n7437);
   U24314 : OAI22_X1 port map( A1 => n30877, A2 => n25445, B1 => n30959, B2 => 
                           n30869, ZN => n7438);
   U24315 : OAI22_X1 port map( A1 => n30877, A2 => n25444, B1 => n30962, B2 => 
                           n30869, ZN => n7439);
   U24316 : OAI22_X1 port map( A1 => n30877, A2 => n25443, B1 => n30965, B2 => 
                           n30869, ZN => n7440);
   U24317 : OAI22_X1 port map( A1 => n30877, A2 => n25442, B1 => n30968, B2 => 
                           n30869, ZN => n7441);
   U24318 : OAI22_X1 port map( A1 => n30877, A2 => n25441, B1 => n30971, B2 => 
                           n30869, ZN => n7442);
   U24319 : OAI22_X1 port map( A1 => n30877, A2 => n25440, B1 => n30974, B2 => 
                           n30869, ZN => n7443);
   U24320 : OAI22_X1 port map( A1 => n30877, A2 => n25439, B1 => n30977, B2 => 
                           n30869, ZN => n7444);
   U24321 : OAI22_X1 port map( A1 => n30878, A2 => n25438, B1 => n30980, B2 => 
                           n30870, ZN => n7445);
   U24322 : OAI22_X1 port map( A1 => n30878, A2 => n25437, B1 => n30983, B2 => 
                           n30870, ZN => n7446);
   U24323 : OAI22_X1 port map( A1 => n30878, A2 => n25436, B1 => n30986, B2 => 
                           n30870, ZN => n7447);
   U24324 : OAI22_X1 port map( A1 => n30878, A2 => n25435, B1 => n30989, B2 => 
                           n30870, ZN => n7448);
   U24325 : OAI22_X1 port map( A1 => n30878, A2 => n25434, B1 => n30992, B2 => 
                           n30870, ZN => n7449);
   U24326 : OAI22_X1 port map( A1 => n30878, A2 => n25433, B1 => n30995, B2 => 
                           n30870, ZN => n7450);
   U24327 : OAI22_X1 port map( A1 => n30878, A2 => n25432, B1 => n30998, B2 => 
                           n30870, ZN => n7451);
   U24328 : OAI22_X1 port map( A1 => n30878, A2 => n25431, B1 => n31001, B2 => 
                           n30870, ZN => n7452);
   U24329 : OAI22_X1 port map( A1 => n30878, A2 => n25430, B1 => n31004, B2 => 
                           n30870, ZN => n7453);
   U24330 : OAI22_X1 port map( A1 => n30878, A2 => n25429, B1 => n31007, B2 => 
                           n30870, ZN => n7454);
   U24331 : OAI22_X1 port map( A1 => n30878, A2 => n25428, B1 => n31010, B2 => 
                           n30870, ZN => n7455);
   U24332 : OAI22_X1 port map( A1 => n30878, A2 => n25427, B1 => n31013, B2 => 
                           n30870, ZN => n7456);
   U24333 : OAI22_X1 port map( A1 => n30878, A2 => n25426, B1 => n31016, B2 => 
                           n30871, ZN => n7457);
   U24334 : OAI22_X1 port map( A1 => n30879, A2 => n25425, B1 => n31019, B2 => 
                           n30871, ZN => n7458);
   U24335 : OAI22_X1 port map( A1 => n30879, A2 => n25424, B1 => n31022, B2 => 
                           n30871, ZN => n7459);
   U24336 : OAI22_X1 port map( A1 => n30879, A2 => n25423, B1 => n31025, B2 => 
                           n30871, ZN => n7460);
   U24337 : OAI22_X1 port map( A1 => n30879, A2 => n25422, B1 => n31028, B2 => 
                           n30871, ZN => n7461);
   U24338 : OAI22_X1 port map( A1 => n30879, A2 => n25421, B1 => n31031, B2 => 
                           n30871, ZN => n7462);
   U24339 : OAI22_X1 port map( A1 => n30879, A2 => n25420, B1 => n31034, B2 => 
                           n30871, ZN => n7463);
   U24340 : OAI22_X1 port map( A1 => n30879, A2 => n25419, B1 => n31037, B2 => 
                           n30871, ZN => n7464);
   U24341 : OAI22_X1 port map( A1 => n30879, A2 => n25418, B1 => n31040, B2 => 
                           n30871, ZN => n7465);
   U24342 : OAI22_X1 port map( A1 => n30879, A2 => n25417, B1 => n31043, B2 => 
                           n30871, ZN => n7466);
   U24343 : OAI22_X1 port map( A1 => n30879, A2 => n25416, B1 => n31046, B2 => 
                           n30871, ZN => n7467);
   U24344 : OAI22_X1 port map( A1 => n30879, A2 => n25415, B1 => n31049, B2 => 
                           n30871, ZN => n7468);
   U24345 : OAI22_X1 port map( A1 => n30879, A2 => n25414, B1 => n31052, B2 => 
                           n30872, ZN => n7469);
   U24346 : OAI22_X1 port map( A1 => n30879, A2 => n25413, B1 => n31055, B2 => 
                           n30872, ZN => n7470);
   U24347 : OAI22_X1 port map( A1 => n30880, A2 => n25412, B1 => n31058, B2 => 
                           n30872, ZN => n7471);
   U24348 : OAI22_X1 port map( A1 => n30880, A2 => n25411, B1 => n31061, B2 => 
                           n30872, ZN => n7472);
   U24349 : OAI22_X1 port map( A1 => n30880, A2 => n25410, B1 => n31064, B2 => 
                           n30872, ZN => n7473);
   U24350 : OAI22_X1 port map( A1 => n30880, A2 => n25409, B1 => n31067, B2 => 
                           n30872, ZN => n7474);
   U24351 : OAI22_X1 port map( A1 => n30880, A2 => n25408, B1 => n31070, B2 => 
                           n30872, ZN => n7475);
   U24352 : OAI22_X1 port map( A1 => n30880, A2 => n25407, B1 => n31073, B2 => 
                           n30872, ZN => n7476);
   U24353 : OAI22_X1 port map( A1 => n30880, A2 => n25406, B1 => n31076, B2 => 
                           n30872, ZN => n7477);
   U24354 : OAI22_X1 port map( A1 => n30880, A2 => n25405, B1 => n31079, B2 => 
                           n30872, ZN => n7478);
   U24355 : OAI22_X1 port map( A1 => n30880, A2 => n25404, B1 => n31082, B2 => 
                           n30872, ZN => n7479);
   U24356 : OAI22_X1 port map( A1 => n30880, A2 => n25403, B1 => n31085, B2 => 
                           n30872, ZN => n7480);
   U24357 : OAI22_X1 port map( A1 => n30880, A2 => n25402, B1 => n31088, B2 => 
                           n30873, ZN => n7481);
   U24358 : OAI22_X1 port map( A1 => n30880, A2 => n25401, B1 => n31091, B2 => 
                           n30873, ZN => n7482);
   U24359 : OAI22_X1 port map( A1 => n30880, A2 => n25400, B1 => n31094, B2 => 
                           n30873, ZN => n7483);
   U24360 : OAI22_X1 port map( A1 => n30881, A2 => n25399, B1 => n31097, B2 => 
                           n30873, ZN => n7484);
   U24361 : OAI22_X1 port map( A1 => n30881, A2 => n25398, B1 => n31100, B2 => 
                           n30873, ZN => n7485);
   U24362 : OAI22_X1 port map( A1 => n30881, A2 => n25397, B1 => n31103, B2 => 
                           n30873, ZN => n7486);
   U24363 : OAI22_X1 port map( A1 => n30881, A2 => n25396, B1 => n31106, B2 => 
                           n30873, ZN => n7487);
   U24364 : OAI22_X1 port map( A1 => n30881, A2 => n25395, B1 => n31109, B2 => 
                           n30873, ZN => n7488);
   U24365 : OAI22_X1 port map( A1 => n30881, A2 => n25394, B1 => n31112, B2 => 
                           n30873, ZN => n7489);
   U24366 : OAI22_X1 port map( A1 => n30881, A2 => n25393, B1 => n31115, B2 => 
                           n30873, ZN => n7490);
   U24367 : OAI22_X1 port map( A1 => n30881, A2 => n25392, B1 => n31118, B2 => 
                           n30873, ZN => n7491);
   U24368 : OAI22_X1 port map( A1 => n30881, A2 => n25391, B1 => n31121, B2 => 
                           n30873, ZN => n7492);
   U24369 : OAI22_X1 port map( A1 => n30752, A2 => n25860, B1 => n30981, B2 => 
                           n30744, ZN => n6805);
   U24370 : OAI22_X1 port map( A1 => n30752, A2 => n25859, B1 => n30984, B2 => 
                           n30744, ZN => n6806);
   U24371 : OAI22_X1 port map( A1 => n30752, A2 => n25858, B1 => n30987, B2 => 
                           n30744, ZN => n6807);
   U24372 : OAI22_X1 port map( A1 => n30752, A2 => n25857, B1 => n30990, B2 => 
                           n30744, ZN => n6808);
   U24373 : OAI22_X1 port map( A1 => n30752, A2 => n25856, B1 => n30993, B2 => 
                           n30744, ZN => n6809);
   U24374 : OAI22_X1 port map( A1 => n30752, A2 => n25855, B1 => n30996, B2 => 
                           n30744, ZN => n6810);
   U24375 : OAI22_X1 port map( A1 => n30752, A2 => n25854, B1 => n30999, B2 => 
                           n30744, ZN => n6811);
   U24376 : OAI22_X1 port map( A1 => n30752, A2 => n25853, B1 => n31002, B2 => 
                           n30744, ZN => n6812);
   U24377 : OAI22_X1 port map( A1 => n30752, A2 => n25852, B1 => n31005, B2 => 
                           n30744, ZN => n6813);
   U24378 : OAI22_X1 port map( A1 => n30752, A2 => n25851, B1 => n31008, B2 => 
                           n30744, ZN => n6814);
   U24379 : OAI22_X1 port map( A1 => n30752, A2 => n25850, B1 => n31011, B2 => 
                           n30744, ZN => n6815);
   U24380 : OAI22_X1 port map( A1 => n30752, A2 => n25849, B1 => n31014, B2 => 
                           n30744, ZN => n6816);
   U24381 : OAI22_X1 port map( A1 => n30752, A2 => n25848, B1 => n31017, B2 => 
                           n30745, ZN => n6817);
   U24382 : OAI22_X1 port map( A1 => n30753, A2 => n25847, B1 => n31020, B2 => 
                           n30745, ZN => n6818);
   U24383 : OAI22_X1 port map( A1 => n30753, A2 => n25846, B1 => n31023, B2 => 
                           n30745, ZN => n6819);
   U24384 : OAI22_X1 port map( A1 => n30753, A2 => n25845, B1 => n31026, B2 => 
                           n30745, ZN => n6820);
   U24385 : OAI22_X1 port map( A1 => n30753, A2 => n25844, B1 => n31029, B2 => 
                           n30745, ZN => n6821);
   U24386 : OAI22_X1 port map( A1 => n30753, A2 => n25843, B1 => n31032, B2 => 
                           n30745, ZN => n6822);
   U24387 : OAI22_X1 port map( A1 => n30753, A2 => n25842, B1 => n31035, B2 => 
                           n30745, ZN => n6823);
   U24388 : OAI22_X1 port map( A1 => n30753, A2 => n25841, B1 => n31038, B2 => 
                           n30745, ZN => n6824);
   U24389 : OAI22_X1 port map( A1 => n30753, A2 => n25840, B1 => n31041, B2 => 
                           n30745, ZN => n6825);
   U24390 : OAI22_X1 port map( A1 => n30753, A2 => n25839, B1 => n31044, B2 => 
                           n30745, ZN => n6826);
   U24391 : OAI22_X1 port map( A1 => n30753, A2 => n25838, B1 => n31047, B2 => 
                           n30745, ZN => n6827);
   U24392 : OAI22_X1 port map( A1 => n30753, A2 => n25837, B1 => n31050, B2 => 
                           n30745, ZN => n6828);
   U24393 : OAI22_X1 port map( A1 => n30753, A2 => n25836, B1 => n31053, B2 => 
                           n30746, ZN => n6829);
   U24394 : OAI22_X1 port map( A1 => n30753, A2 => n25835, B1 => n31056, B2 => 
                           n30746, ZN => n6830);
   U24395 : OAI22_X1 port map( A1 => n30754, A2 => n25834, B1 => n31059, B2 => 
                           n30746, ZN => n6831);
   U24396 : OAI22_X1 port map( A1 => n30754, A2 => n25833, B1 => n31062, B2 => 
                           n30746, ZN => n6832);
   U24397 : OAI22_X1 port map( A1 => n30754, A2 => n25832, B1 => n31065, B2 => 
                           n30746, ZN => n6833);
   U24398 : OAI22_X1 port map( A1 => n30754, A2 => n25831, B1 => n31068, B2 => 
                           n30746, ZN => n6834);
   U24399 : OAI22_X1 port map( A1 => n30754, A2 => n25830, B1 => n31071, B2 => 
                           n30746, ZN => n6835);
   U24400 : OAI22_X1 port map( A1 => n30754, A2 => n25829, B1 => n31074, B2 => 
                           n30746, ZN => n6836);
   U24401 : OAI22_X1 port map( A1 => n30754, A2 => n25828, B1 => n31077, B2 => 
                           n30746, ZN => n6837);
   U24402 : OAI22_X1 port map( A1 => n30754, A2 => n25827, B1 => n31080, B2 => 
                           n30746, ZN => n6838);
   U24403 : OAI22_X1 port map( A1 => n30754, A2 => n25826, B1 => n31083, B2 => 
                           n30746, ZN => n6839);
   U24404 : OAI22_X1 port map( A1 => n30754, A2 => n25825, B1 => n31086, B2 => 
                           n30746, ZN => n6840);
   U24405 : OAI22_X1 port map( A1 => n30754, A2 => n25824, B1 => n31089, B2 => 
                           n30747, ZN => n6841);
   U24406 : OAI22_X1 port map( A1 => n30754, A2 => n25823, B1 => n31092, B2 => 
                           n30747, ZN => n6842);
   U24407 : OAI22_X1 port map( A1 => n30754, A2 => n25822, B1 => n31095, B2 => 
                           n30747, ZN => n6843);
   U24408 : OAI22_X1 port map( A1 => n30755, A2 => n25821, B1 => n31098, B2 => 
                           n30747, ZN => n6844);
   U24409 : OAI22_X1 port map( A1 => n30755, A2 => n25820, B1 => n31101, B2 => 
                           n30747, ZN => n6845);
   U24410 : OAI22_X1 port map( A1 => n30755, A2 => n25819, B1 => n31104, B2 => 
                           n30747, ZN => n6846);
   U24411 : OAI22_X1 port map( A1 => n30755, A2 => n25818, B1 => n31107, B2 => 
                           n30747, ZN => n6847);
   U24412 : OAI22_X1 port map( A1 => n30755, A2 => n25817, B1 => n31110, B2 => 
                           n30747, ZN => n6848);
   U24413 : OAI22_X1 port map( A1 => n30755, A2 => n25816, B1 => n31113, B2 => 
                           n30747, ZN => n6849);
   U24414 : OAI22_X1 port map( A1 => n30755, A2 => n25815, B1 => n31116, B2 => 
                           n30747, ZN => n6850);
   U24415 : OAI22_X1 port map( A1 => n30755, A2 => n25814, B1 => n31119, B2 => 
                           n30747, ZN => n6851);
   U24416 : OAI22_X1 port map( A1 => n30755, A2 => n25813, B1 => n31122, B2 => 
                           n30747, ZN => n6852);
   U24417 : OAI22_X1 port map( A1 => n30751, A2 => n25872, B1 => n30945, B2 => 
                           n30743, ZN => n6793);
   U24418 : OAI22_X1 port map( A1 => n30751, A2 => n25871, B1 => n30948, B2 => 
                           n30743, ZN => n6794);
   U24419 : OAI22_X1 port map( A1 => n30751, A2 => n25870, B1 => n30951, B2 => 
                           n30743, ZN => n6795);
   U24420 : OAI22_X1 port map( A1 => n30751, A2 => n25869, B1 => n30954, B2 => 
                           n30743, ZN => n6796);
   U24421 : OAI22_X1 port map( A1 => n30751, A2 => n25868, B1 => n30957, B2 => 
                           n30743, ZN => n6797);
   U24422 : OAI22_X1 port map( A1 => n30751, A2 => n25867, B1 => n30960, B2 => 
                           n30743, ZN => n6798);
   U24423 : OAI22_X1 port map( A1 => n30751, A2 => n25866, B1 => n30963, B2 => 
                           n30743, ZN => n6799);
   U24424 : OAI22_X1 port map( A1 => n30751, A2 => n25865, B1 => n30966, B2 => 
                           n30743, ZN => n6800);
   U24425 : OAI22_X1 port map( A1 => n30751, A2 => n25864, B1 => n30969, B2 => 
                           n30743, ZN => n6801);
   U24426 : OAI22_X1 port map( A1 => n30751, A2 => n25863, B1 => n30972, B2 => 
                           n30743, ZN => n6802);
   U24427 : OAI22_X1 port map( A1 => n30751, A2 => n25862, B1 => n30975, B2 => 
                           n30743, ZN => n6803);
   U24428 : OAI22_X1 port map( A1 => n30751, A2 => n25861, B1 => n30978, B2 => 
                           n30743, ZN => n6804);
   U24429 : OAI22_X1 port map( A1 => n18111, A2 => n30675, B1 => n30981, B2 => 
                           n30669, ZN => n6421);
   U24430 : OAI22_X1 port map( A1 => n18110, A2 => n30675, B1 => n30984, B2 => 
                           n30669, ZN => n6422);
   U24431 : OAI22_X1 port map( A1 => n18109, A2 => n30675, B1 => n30987, B2 => 
                           n30669, ZN => n6423);
   U24432 : OAI22_X1 port map( A1 => n18108, A2 => n30675, B1 => n30990, B2 => 
                           n30669, ZN => n6424);
   U24433 : OAI22_X1 port map( A1 => n18107, A2 => n30675, B1 => n30993, B2 => 
                           n30669, ZN => n6425);
   U24434 : OAI22_X1 port map( A1 => n18106, A2 => n30675, B1 => n30996, B2 => 
                           n30669, ZN => n6426);
   U24435 : OAI22_X1 port map( A1 => n18105, A2 => n30675, B1 => n30999, B2 => 
                           n30669, ZN => n6427);
   U24436 : OAI22_X1 port map( A1 => n18104, A2 => n30675, B1 => n31002, B2 => 
                           n30669, ZN => n6428);
   U24437 : OAI22_X1 port map( A1 => n18103, A2 => n30675, B1 => n31005, B2 => 
                           n30669, ZN => n6429);
   U24438 : OAI22_X1 port map( A1 => n18102, A2 => n30675, B1 => n31008, B2 => 
                           n30669, ZN => n6430);
   U24439 : OAI22_X1 port map( A1 => n18101, A2 => n30675, B1 => n31011, B2 => 
                           n30669, ZN => n6431);
   U24440 : OAI22_X1 port map( A1 => n18100, A2 => n30676, B1 => n31014, B2 => 
                           n30669, ZN => n6432);
   U24441 : OAI22_X1 port map( A1 => n18099, A2 => n30676, B1 => n31017, B2 => 
                           n30670, ZN => n6433);
   U24442 : OAI22_X1 port map( A1 => n18098, A2 => n30676, B1 => n31020, B2 => 
                           n30670, ZN => n6434);
   U24443 : OAI22_X1 port map( A1 => n18097, A2 => n30676, B1 => n31023, B2 => 
                           n30670, ZN => n6435);
   U24444 : OAI22_X1 port map( A1 => n18096, A2 => n30676, B1 => n31026, B2 => 
                           n30670, ZN => n6436);
   U24445 : OAI22_X1 port map( A1 => n18095, A2 => n30676, B1 => n31029, B2 => 
                           n30670, ZN => n6437);
   U24446 : OAI22_X1 port map( A1 => n18094, A2 => n30676, B1 => n31032, B2 => 
                           n30670, ZN => n6438);
   U24447 : OAI22_X1 port map( A1 => n18093, A2 => n30676, B1 => n31035, B2 => 
                           n30670, ZN => n6439);
   U24448 : OAI22_X1 port map( A1 => n18092, A2 => n30676, B1 => n31038, B2 => 
                           n30670, ZN => n6440);
   U24449 : OAI22_X1 port map( A1 => n18091, A2 => n30676, B1 => n31041, B2 => 
                           n30670, ZN => n6441);
   U24450 : OAI22_X1 port map( A1 => n18090, A2 => n30676, B1 => n31044, B2 => 
                           n30670, ZN => n6442);
   U24451 : OAI22_X1 port map( A1 => n18089, A2 => n30676, B1 => n31047, B2 => 
                           n30670, ZN => n6443);
   U24452 : OAI22_X1 port map( A1 => n18088, A2 => n30677, B1 => n31050, B2 => 
                           n30670, ZN => n6444);
   U24453 : OAI22_X1 port map( A1 => n18087, A2 => n30677, B1 => n31053, B2 => 
                           n30671, ZN => n6445);
   U24454 : OAI22_X1 port map( A1 => n18086, A2 => n30677, B1 => n31056, B2 => 
                           n30671, ZN => n6446);
   U24455 : OAI22_X1 port map( A1 => n18085, A2 => n30677, B1 => n31059, B2 => 
                           n30671, ZN => n6447);
   U24456 : OAI22_X1 port map( A1 => n18084, A2 => n30677, B1 => n31062, B2 => 
                           n30671, ZN => n6448);
   U24457 : OAI22_X1 port map( A1 => n18083, A2 => n30677, B1 => n31065, B2 => 
                           n30671, ZN => n6449);
   U24458 : OAI22_X1 port map( A1 => n18082, A2 => n30677, B1 => n31068, B2 => 
                           n30671, ZN => n6450);
   U24459 : OAI22_X1 port map( A1 => n18081, A2 => n30677, B1 => n31071, B2 => 
                           n30671, ZN => n6451);
   U24460 : OAI22_X1 port map( A1 => n18080, A2 => n30677, B1 => n31074, B2 => 
                           n30671, ZN => n6452);
   U24461 : OAI22_X1 port map( A1 => n18079, A2 => n30677, B1 => n31077, B2 => 
                           n30671, ZN => n6453);
   U24462 : OAI22_X1 port map( A1 => n18078, A2 => n30677, B1 => n31080, B2 => 
                           n30671, ZN => n6454);
   U24463 : OAI22_X1 port map( A1 => n18077, A2 => n30677, B1 => n31083, B2 => 
                           n30671, ZN => n6455);
   U24464 : OAI22_X1 port map( A1 => n18076, A2 => n30678, B1 => n31086, B2 => 
                           n30671, ZN => n6456);
   U24465 : OAI22_X1 port map( A1 => n18075, A2 => n30678, B1 => n31089, B2 => 
                           n30672, ZN => n6457);
   U24466 : OAI22_X1 port map( A1 => n18074, A2 => n30678, B1 => n31092, B2 => 
                           n30672, ZN => n6458);
   U24467 : OAI22_X1 port map( A1 => n18073, A2 => n30678, B1 => n31095, B2 => 
                           n30672, ZN => n6459);
   U24468 : OAI22_X1 port map( A1 => n18072, A2 => n30678, B1 => n31098, B2 => 
                           n30672, ZN => n6460);
   U24469 : OAI22_X1 port map( A1 => n18071, A2 => n30678, B1 => n31101, B2 => 
                           n30672, ZN => n6461);
   U24470 : OAI22_X1 port map( A1 => n18070, A2 => n30678, B1 => n31104, B2 => 
                           n30672, ZN => n6462);
   U24471 : OAI22_X1 port map( A1 => n18069, A2 => n30678, B1 => n31107, B2 => 
                           n30672, ZN => n6463);
   U24472 : OAI22_X1 port map( A1 => n18068, A2 => n30678, B1 => n31110, B2 => 
                           n30672, ZN => n6464);
   U24473 : OAI22_X1 port map( A1 => n18067, A2 => n30678, B1 => n31113, B2 => 
                           n30672, ZN => n6465);
   U24474 : OAI22_X1 port map( A1 => n18066, A2 => n30678, B1 => n31116, B2 => 
                           n30672, ZN => n6466);
   U24475 : OAI22_X1 port map( A1 => n18065, A2 => n30678, B1 => n31119, B2 => 
                           n30672, ZN => n6467);
   U24476 : OAI22_X1 port map( A1 => n18064, A2 => n30679, B1 => n31122, B2 => 
                           n30672, ZN => n6468);
   U24477 : OAI22_X1 port map( A1 => n18123, A2 => n30674, B1 => n30945, B2 => 
                           n30668, ZN => n6409);
   U24478 : OAI22_X1 port map( A1 => n18122, A2 => n30674, B1 => n30948, B2 => 
                           n30668, ZN => n6410);
   U24479 : OAI22_X1 port map( A1 => n18121, A2 => n30674, B1 => n30951, B2 => 
                           n30668, ZN => n6411);
   U24480 : OAI22_X1 port map( A1 => n18120, A2 => n30674, B1 => n30954, B2 => 
                           n30668, ZN => n6412);
   U24481 : OAI22_X1 port map( A1 => n18119, A2 => n30674, B1 => n30957, B2 => 
                           n30668, ZN => n6413);
   U24482 : OAI22_X1 port map( A1 => n18118, A2 => n30674, B1 => n30960, B2 => 
                           n30668, ZN => n6414);
   U24483 : OAI22_X1 port map( A1 => n18117, A2 => n30674, B1 => n30963, B2 => 
                           n30668, ZN => n6415);
   U24484 : OAI22_X1 port map( A1 => n18116, A2 => n30674, B1 => n30966, B2 => 
                           n30668, ZN => n6416);
   U24485 : OAI22_X1 port map( A1 => n18115, A2 => n30674, B1 => n30969, B2 => 
                           n30668, ZN => n6417);
   U24486 : OAI22_X1 port map( A1 => n18114, A2 => n30674, B1 => n30972, B2 => 
                           n30668, ZN => n6418);
   U24487 : OAI22_X1 port map( A1 => n18113, A2 => n30674, B1 => n30975, B2 => 
                           n30668, ZN => n6419);
   U24488 : OAI22_X1 port map( A1 => n18112, A2 => n30675, B1 => n30978, B2 => 
                           n30668, ZN => n6420);
   U24489 : OAI22_X1 port map( A1 => n9288, A2 => n30712, B1 => n30945, B2 => 
                           n30706, ZN => n6601);
   U24490 : OAI22_X1 port map( A1 => n9283, A2 => n30712, B1 => n30948, B2 => 
                           n30706, ZN => n6602);
   U24491 : OAI22_X1 port map( A1 => n9278, A2 => n30712, B1 => n30951, B2 => 
                           n30706, ZN => n6603);
   U24492 : OAI22_X1 port map( A1 => n9273, A2 => n30712, B1 => n30954, B2 => 
                           n30706, ZN => n6604);
   U24493 : OAI22_X1 port map( A1 => n9268, A2 => n30712, B1 => n30957, B2 => 
                           n30706, ZN => n6605);
   U24494 : OAI22_X1 port map( A1 => n9263, A2 => n30712, B1 => n30960, B2 => 
                           n30706, ZN => n6606);
   U24495 : OAI22_X1 port map( A1 => n9258, A2 => n30712, B1 => n30963, B2 => 
                           n30706, ZN => n6607);
   U24496 : OAI22_X1 port map( A1 => n9253, A2 => n30712, B1 => n30966, B2 => 
                           n30706, ZN => n6608);
   U24497 : OAI22_X1 port map( A1 => n9248, A2 => n30712, B1 => n30969, B2 => 
                           n30706, ZN => n6609);
   U24498 : OAI22_X1 port map( A1 => n9243, A2 => n30712, B1 => n30972, B2 => 
                           n30706, ZN => n6610);
   U24499 : OAI22_X1 port map( A1 => n9238, A2 => n30712, B1 => n30975, B2 => 
                           n30706, ZN => n6611);
   U24500 : OAI22_X1 port map( A1 => n9233, A2 => n30713, B1 => n30978, B2 => 
                           n30706, ZN => n6612);
   U24501 : OAI22_X1 port map( A1 => n9228, A2 => n30713, B1 => n30981, B2 => 
                           n30707, ZN => n6613);
   U24502 : OAI22_X1 port map( A1 => n9223, A2 => n30713, B1 => n30984, B2 => 
                           n30707, ZN => n6614);
   U24503 : OAI22_X1 port map( A1 => n9218, A2 => n30713, B1 => n30987, B2 => 
                           n30707, ZN => n6615);
   U24504 : OAI22_X1 port map( A1 => n9213, A2 => n30713, B1 => n30990, B2 => 
                           n30707, ZN => n6616);
   U24505 : OAI22_X1 port map( A1 => n9208, A2 => n30713, B1 => n30993, B2 => 
                           n30707, ZN => n6617);
   U24506 : OAI22_X1 port map( A1 => n9203, A2 => n30713, B1 => n30996, B2 => 
                           n30707, ZN => n6618);
   U24507 : OAI22_X1 port map( A1 => n9198, A2 => n30713, B1 => n30999, B2 => 
                           n30707, ZN => n6619);
   U24508 : OAI22_X1 port map( A1 => n9193, A2 => n30713, B1 => n31002, B2 => 
                           n30707, ZN => n6620);
   U24509 : OAI22_X1 port map( A1 => n9188, A2 => n30713, B1 => n31005, B2 => 
                           n30707, ZN => n6621);
   U24510 : OAI22_X1 port map( A1 => n9183, A2 => n30713, B1 => n31008, B2 => 
                           n30707, ZN => n6622);
   U24511 : OAI22_X1 port map( A1 => n9178, A2 => n30713, B1 => n31011, B2 => 
                           n30707, ZN => n6623);
   U24512 : OAI22_X1 port map( A1 => n9173, A2 => n30714, B1 => n31014, B2 => 
                           n30707, ZN => n6624);
   U24513 : OAI22_X1 port map( A1 => n9168, A2 => n30714, B1 => n31017, B2 => 
                           n30708, ZN => n6625);
   U24514 : OAI22_X1 port map( A1 => n9163, A2 => n30714, B1 => n31020, B2 => 
                           n30708, ZN => n6626);
   U24515 : OAI22_X1 port map( A1 => n9158, A2 => n30714, B1 => n31023, B2 => 
                           n30708, ZN => n6627);
   U24516 : OAI22_X1 port map( A1 => n9153, A2 => n30714, B1 => n31026, B2 => 
                           n30708, ZN => n6628);
   U24517 : OAI22_X1 port map( A1 => n9148, A2 => n30714, B1 => n31029, B2 => 
                           n30708, ZN => n6629);
   U24518 : OAI22_X1 port map( A1 => n9143, A2 => n30714, B1 => n31032, B2 => 
                           n30708, ZN => n6630);
   U24519 : OAI22_X1 port map( A1 => n9138, A2 => n30714, B1 => n31035, B2 => 
                           n30708, ZN => n6631);
   U24520 : OAI22_X1 port map( A1 => n9133, A2 => n30714, B1 => n31038, B2 => 
                           n30708, ZN => n6632);
   U24521 : OAI22_X1 port map( A1 => n9128, A2 => n30714, B1 => n31041, B2 => 
                           n30708, ZN => n6633);
   U24522 : OAI22_X1 port map( A1 => n9123, A2 => n30714, B1 => n31044, B2 => 
                           n30708, ZN => n6634);
   U24523 : OAI22_X1 port map( A1 => n9118, A2 => n30714, B1 => n31047, B2 => 
                           n30708, ZN => n6635);
   U24524 : OAI22_X1 port map( A1 => n9113, A2 => n30715, B1 => n31050, B2 => 
                           n30708, ZN => n6636);
   U24525 : OAI22_X1 port map( A1 => n9108, A2 => n30715, B1 => n31053, B2 => 
                           n30709, ZN => n6637);
   U24526 : OAI22_X1 port map( A1 => n9103, A2 => n30715, B1 => n31056, B2 => 
                           n30709, ZN => n6638);
   U24527 : OAI22_X1 port map( A1 => n9098, A2 => n30715, B1 => n31059, B2 => 
                           n30709, ZN => n6639);
   U24528 : OAI22_X1 port map( A1 => n9093, A2 => n30715, B1 => n31062, B2 => 
                           n30709, ZN => n6640);
   U24529 : OAI22_X1 port map( A1 => n9088, A2 => n30715, B1 => n31065, B2 => 
                           n30709, ZN => n6641);
   U24530 : OAI22_X1 port map( A1 => n9083, A2 => n30715, B1 => n31068, B2 => 
                           n30709, ZN => n6642);
   U24531 : OAI22_X1 port map( A1 => n9078, A2 => n30715, B1 => n31071, B2 => 
                           n30709, ZN => n6643);
   U24532 : OAI22_X1 port map( A1 => n9073, A2 => n30715, B1 => n31074, B2 => 
                           n30709, ZN => n6644);
   U24533 : OAI22_X1 port map( A1 => n9068, A2 => n30715, B1 => n31077, B2 => 
                           n30709, ZN => n6645);
   U24534 : OAI22_X1 port map( A1 => n9063, A2 => n30715, B1 => n31080, B2 => 
                           n30709, ZN => n6646);
   U24535 : OAI22_X1 port map( A1 => n9058, A2 => n30715, B1 => n31083, B2 => 
                           n30709, ZN => n6647);
   U24536 : OAI22_X1 port map( A1 => n9053, A2 => n30716, B1 => n31086, B2 => 
                           n30709, ZN => n6648);
   U24537 : OAI22_X1 port map( A1 => n9048, A2 => n30716, B1 => n31089, B2 => 
                           n30710, ZN => n6649);
   U24538 : OAI22_X1 port map( A1 => n9043, A2 => n30716, B1 => n31092, B2 => 
                           n30710, ZN => n6650);
   U24539 : OAI22_X1 port map( A1 => n9038, A2 => n30716, B1 => n31095, B2 => 
                           n30710, ZN => n6651);
   U24540 : OAI22_X1 port map( A1 => n9033, A2 => n30716, B1 => n31098, B2 => 
                           n30710, ZN => n6652);
   U24541 : OAI22_X1 port map( A1 => n9028, A2 => n30716, B1 => n31101, B2 => 
                           n30710, ZN => n6653);
   U24542 : OAI22_X1 port map( A1 => n9023, A2 => n30716, B1 => n31104, B2 => 
                           n30710, ZN => n6654);
   U24543 : OAI22_X1 port map( A1 => n9018, A2 => n30716, B1 => n31107, B2 => 
                           n30710, ZN => n6655);
   U24544 : OAI22_X1 port map( A1 => n9013, A2 => n30716, B1 => n31110, B2 => 
                           n30710, ZN => n6656);
   U24545 : OAI22_X1 port map( A1 => n9008, A2 => n30716, B1 => n31113, B2 => 
                           n30710, ZN => n6657);
   U24546 : OAI22_X1 port map( A1 => n9003, A2 => n30716, B1 => n31116, B2 => 
                           n30710, ZN => n6658);
   U24547 : OAI22_X1 port map( A1 => n8998, A2 => n30716, B1 => n31119, B2 => 
                           n30710, ZN => n6659);
   U24548 : OAI22_X1 port map( A1 => n8993, A2 => n30717, B1 => n31122, B2 => 
                           n30710, ZN => n6660);
   U24549 : OAI22_X1 port map( A1 => n9996, A2 => n30728, B1 => n30981, B2 => 
                           n30719, ZN => n6677);
   U24550 : OAI22_X1 port map( A1 => n9991, A2 => n30728, B1 => n30984, B2 => 
                           n30719, ZN => n6678);
   U24551 : OAI22_X1 port map( A1 => n9986, A2 => n30728, B1 => n30987, B2 => 
                           n30719, ZN => n6679);
   U24552 : OAI22_X1 port map( A1 => n9981, A2 => n30728, B1 => n30990, B2 => 
                           n30719, ZN => n6680);
   U24553 : OAI22_X1 port map( A1 => n9976, A2 => n30728, B1 => n30993, B2 => 
                           n30719, ZN => n6681);
   U24554 : OAI22_X1 port map( A1 => n9971, A2 => n30727, B1 => n30996, B2 => 
                           n30719, ZN => n6682);
   U24555 : OAI22_X1 port map( A1 => n9966, A2 => n30727, B1 => n30999, B2 => 
                           n30719, ZN => n6683);
   U24556 : OAI22_X1 port map( A1 => n9961, A2 => n30727, B1 => n31002, B2 => 
                           n30719, ZN => n6684);
   U24557 : OAI22_X1 port map( A1 => n9956, A2 => n30727, B1 => n31005, B2 => 
                           n30719, ZN => n6685);
   U24558 : OAI22_X1 port map( A1 => n9951, A2 => n30727, B1 => n31008, B2 => 
                           n30719, ZN => n6686);
   U24559 : OAI22_X1 port map( A1 => n9946, A2 => n30727, B1 => n31011, B2 => 
                           n30719, ZN => n6687);
   U24560 : OAI22_X1 port map( A1 => n9941, A2 => n30727, B1 => n31014, B2 => 
                           n30719, ZN => n6688);
   U24561 : OAI22_X1 port map( A1 => n9936, A2 => n30727, B1 => n31017, B2 => 
                           n30720, ZN => n6689);
   U24562 : OAI22_X1 port map( A1 => n9931, A2 => n30727, B1 => n31020, B2 => 
                           n30720, ZN => n6690);
   U24563 : OAI22_X1 port map( A1 => n9926, A2 => n30727, B1 => n31023, B2 => 
                           n30720, ZN => n6691);
   U24564 : OAI22_X1 port map( A1 => n9921, A2 => n30727, B1 => n31026, B2 => 
                           n30720, ZN => n6692);
   U24565 : OAI22_X1 port map( A1 => n9916, A2 => n30727, B1 => n31029, B2 => 
                           n30720, ZN => n6693);
   U24566 : OAI22_X1 port map( A1 => n9911, A2 => n30726, B1 => n31032, B2 => 
                           n30720, ZN => n6694);
   U24567 : OAI22_X1 port map( A1 => n9906, A2 => n30726, B1 => n31035, B2 => 
                           n30720, ZN => n6695);
   U24568 : OAI22_X1 port map( A1 => n9901, A2 => n30726, B1 => n31038, B2 => 
                           n30720, ZN => n6696);
   U24569 : OAI22_X1 port map( A1 => n9896, A2 => n30726, B1 => n31041, B2 => 
                           n30720, ZN => n6697);
   U24570 : OAI22_X1 port map( A1 => n9891, A2 => n30726, B1 => n31044, B2 => 
                           n30720, ZN => n6698);
   U24571 : OAI22_X1 port map( A1 => n9886, A2 => n30726, B1 => n31047, B2 => 
                           n30720, ZN => n6699);
   U24572 : OAI22_X1 port map( A1 => n9881, A2 => n30726, B1 => n31050, B2 => 
                           n30720, ZN => n6700);
   U24573 : OAI22_X1 port map( A1 => n9876, A2 => n30726, B1 => n31053, B2 => 
                           n30721, ZN => n6701);
   U24574 : OAI22_X1 port map( A1 => n9871, A2 => n30726, B1 => n31056, B2 => 
                           n30721, ZN => n6702);
   U24575 : OAI22_X1 port map( A1 => n9866, A2 => n30726, B1 => n31059, B2 => 
                           n30721, ZN => n6703);
   U24576 : OAI22_X1 port map( A1 => n9861, A2 => n30726, B1 => n31062, B2 => 
                           n30721, ZN => n6704);
   U24577 : OAI22_X1 port map( A1 => n9856, A2 => n30725, B1 => n31065, B2 => 
                           n30721, ZN => n6705);
   U24578 : OAI22_X1 port map( A1 => n9851, A2 => n30725, B1 => n31068, B2 => 
                           n30721, ZN => n6706);
   U24579 : OAI22_X1 port map( A1 => n9846, A2 => n30725, B1 => n31071, B2 => 
                           n30721, ZN => n6707);
   U24580 : OAI22_X1 port map( A1 => n9841, A2 => n30725, B1 => n31074, B2 => 
                           n30721, ZN => n6708);
   U24581 : OAI22_X1 port map( A1 => n9836, A2 => n30725, B1 => n31077, B2 => 
                           n30721, ZN => n6709);
   U24582 : OAI22_X1 port map( A1 => n9831, A2 => n30725, B1 => n31080, B2 => 
                           n30721, ZN => n6710);
   U24583 : OAI22_X1 port map( A1 => n9826, A2 => n30725, B1 => n31083, B2 => 
                           n30721, ZN => n6711);
   U24584 : OAI22_X1 port map( A1 => n9821, A2 => n30725, B1 => n31086, B2 => 
                           n30721, ZN => n6712);
   U24585 : OAI22_X1 port map( A1 => n9816, A2 => n30725, B1 => n31089, B2 => 
                           n30722, ZN => n6713);
   U24586 : OAI22_X1 port map( A1 => n9811, A2 => n30725, B1 => n31092, B2 => 
                           n30722, ZN => n6714);
   U24587 : OAI22_X1 port map( A1 => n9806, A2 => n30725, B1 => n31095, B2 => 
                           n30722, ZN => n6715);
   U24588 : OAI22_X1 port map( A1 => n9801, A2 => n30725, B1 => n31098, B2 => 
                           n30722, ZN => n6716);
   U24589 : OAI22_X1 port map( A1 => n9796, A2 => n30724, B1 => n31101, B2 => 
                           n30722, ZN => n6717);
   U24590 : OAI22_X1 port map( A1 => n9791, A2 => n30724, B1 => n31104, B2 => 
                           n30722, ZN => n6718);
   U24591 : OAI22_X1 port map( A1 => n9786, A2 => n30724, B1 => n31107, B2 => 
                           n30722, ZN => n6719);
   U24592 : OAI22_X1 port map( A1 => n9781, A2 => n30724, B1 => n31110, B2 => 
                           n30722, ZN => n6720);
   U24593 : OAI22_X1 port map( A1 => n9776, A2 => n30724, B1 => n31113, B2 => 
                           n30722, ZN => n6721);
   U24594 : OAI22_X1 port map( A1 => n9771, A2 => n30724, B1 => n31116, B2 => 
                           n30722, ZN => n6722);
   U24595 : OAI22_X1 port map( A1 => n9766, A2 => n30724, B1 => n31119, B2 => 
                           n30722, ZN => n6723);
   U24596 : OAI22_X1 port map( A1 => n9761, A2 => n30724, B1 => n31122, B2 => 
                           n30722, ZN => n6724);
   U24597 : OAI22_X1 port map( A1 => n30738, A2 => n25939, B1 => n30945, B2 => 
                           n30730, ZN => n6729);
   U24598 : OAI22_X1 port map( A1 => n30738, A2 => n25938, B1 => n30948, B2 => 
                           n30730, ZN => n6730);
   U24599 : OAI22_X1 port map( A1 => n30738, A2 => n25937, B1 => n30951, B2 => 
                           n30730, ZN => n6731);
   U24600 : OAI22_X1 port map( A1 => n30738, A2 => n25936, B1 => n30954, B2 => 
                           n30730, ZN => n6732);
   U24601 : OAI22_X1 port map( A1 => n30738, A2 => n25935, B1 => n30957, B2 => 
                           n30730, ZN => n6733);
   U24602 : OAI22_X1 port map( A1 => n30738, A2 => n25934, B1 => n30960, B2 => 
                           n30730, ZN => n6734);
   U24603 : OAI22_X1 port map( A1 => n30738, A2 => n25933, B1 => n30963, B2 => 
                           n30730, ZN => n6735);
   U24604 : OAI22_X1 port map( A1 => n30738, A2 => n25932, B1 => n30966, B2 => 
                           n30730, ZN => n6736);
   U24605 : OAI22_X1 port map( A1 => n30738, A2 => n25931, B1 => n30969, B2 => 
                           n30730, ZN => n6737);
   U24606 : OAI22_X1 port map( A1 => n30738, A2 => n25930, B1 => n30972, B2 => 
                           n30730, ZN => n6738);
   U24607 : OAI22_X1 port map( A1 => n30738, A2 => n25929, B1 => n30975, B2 => 
                           n30730, ZN => n6739);
   U24608 : OAI22_X1 port map( A1 => n30738, A2 => n25928, B1 => n30978, B2 => 
                           n30730, ZN => n6740);
   U24609 : OAI22_X1 port map( A1 => n30739, A2 => n25927, B1 => n30981, B2 => 
                           n30731, ZN => n6741);
   U24610 : OAI22_X1 port map( A1 => n30739, A2 => n25926, B1 => n30984, B2 => 
                           n30731, ZN => n6742);
   U24611 : OAI22_X1 port map( A1 => n30739, A2 => n25925, B1 => n30987, B2 => 
                           n30731, ZN => n6743);
   U24612 : OAI22_X1 port map( A1 => n30739, A2 => n25924, B1 => n30990, B2 => 
                           n30731, ZN => n6744);
   U24613 : OAI22_X1 port map( A1 => n30739, A2 => n25923, B1 => n30993, B2 => 
                           n30731, ZN => n6745);
   U24614 : OAI22_X1 port map( A1 => n30739, A2 => n25922, B1 => n30996, B2 => 
                           n30731, ZN => n6746);
   U24615 : OAI22_X1 port map( A1 => n30739, A2 => n25921, B1 => n30999, B2 => 
                           n30731, ZN => n6747);
   U24616 : OAI22_X1 port map( A1 => n30739, A2 => n25920, B1 => n31002, B2 => 
                           n30731, ZN => n6748);
   U24617 : OAI22_X1 port map( A1 => n30739, A2 => n25919, B1 => n31005, B2 => 
                           n30731, ZN => n6749);
   U24618 : OAI22_X1 port map( A1 => n30739, A2 => n25918, B1 => n31008, B2 => 
                           n30731, ZN => n6750);
   U24619 : OAI22_X1 port map( A1 => n30739, A2 => n25917, B1 => n31011, B2 => 
                           n30731, ZN => n6751);
   U24620 : OAI22_X1 port map( A1 => n30739, A2 => n25916, B1 => n31014, B2 => 
                           n30731, ZN => n6752);
   U24621 : OAI22_X1 port map( A1 => n30739, A2 => n25915, B1 => n31017, B2 => 
                           n30732, ZN => n6753);
   U24622 : OAI22_X1 port map( A1 => n30740, A2 => n25914, B1 => n31020, B2 => 
                           n30732, ZN => n6754);
   U24623 : OAI22_X1 port map( A1 => n30740, A2 => n25913, B1 => n31023, B2 => 
                           n30732, ZN => n6755);
   U24624 : OAI22_X1 port map( A1 => n30740, A2 => n25912, B1 => n31026, B2 => 
                           n30732, ZN => n6756);
   U24625 : OAI22_X1 port map( A1 => n30740, A2 => n25911, B1 => n31029, B2 => 
                           n30732, ZN => n6757);
   U24626 : OAI22_X1 port map( A1 => n30740, A2 => n25910, B1 => n31032, B2 => 
                           n30732, ZN => n6758);
   U24627 : OAI22_X1 port map( A1 => n30740, A2 => n25909, B1 => n31035, B2 => 
                           n30732, ZN => n6759);
   U24628 : OAI22_X1 port map( A1 => n30740, A2 => n25908, B1 => n31038, B2 => 
                           n30732, ZN => n6760);
   U24629 : OAI22_X1 port map( A1 => n30740, A2 => n25907, B1 => n31041, B2 => 
                           n30732, ZN => n6761);
   U24630 : OAI22_X1 port map( A1 => n30740, A2 => n25906, B1 => n31044, B2 => 
                           n30732, ZN => n6762);
   U24631 : OAI22_X1 port map( A1 => n30740, A2 => n25905, B1 => n31047, B2 => 
                           n30732, ZN => n6763);
   U24632 : OAI22_X1 port map( A1 => n30740, A2 => n25904, B1 => n31050, B2 => 
                           n30732, ZN => n6764);
   U24633 : OAI22_X1 port map( A1 => n30740, A2 => n25903, B1 => n31053, B2 => 
                           n30733, ZN => n6765);
   U24634 : OAI22_X1 port map( A1 => n30740, A2 => n25902, B1 => n31056, B2 => 
                           n30733, ZN => n6766);
   U24635 : OAI22_X1 port map( A1 => n30741, A2 => n25901, B1 => n31059, B2 => 
                           n30733, ZN => n6767);
   U24636 : OAI22_X1 port map( A1 => n30741, A2 => n25900, B1 => n31062, B2 => 
                           n30733, ZN => n6768);
   U24637 : OAI22_X1 port map( A1 => n30741, A2 => n25899, B1 => n31065, B2 => 
                           n30733, ZN => n6769);
   U24638 : OAI22_X1 port map( A1 => n30741, A2 => n25898, B1 => n31068, B2 => 
                           n30733, ZN => n6770);
   U24639 : OAI22_X1 port map( A1 => n30741, A2 => n25897, B1 => n31071, B2 => 
                           n30733, ZN => n6771);
   U24640 : OAI22_X1 port map( A1 => n30741, A2 => n25896, B1 => n31074, B2 => 
                           n30733, ZN => n6772);
   U24641 : OAI22_X1 port map( A1 => n30741, A2 => n25895, B1 => n31077, B2 => 
                           n30733, ZN => n6773);
   U24642 : OAI22_X1 port map( A1 => n30741, A2 => n25894, B1 => n31080, B2 => 
                           n30733, ZN => n6774);
   U24643 : OAI22_X1 port map( A1 => n30741, A2 => n25893, B1 => n31083, B2 => 
                           n30733, ZN => n6775);
   U24644 : OAI22_X1 port map( A1 => n30741, A2 => n25892, B1 => n31086, B2 => 
                           n30733, ZN => n6776);
   U24645 : OAI22_X1 port map( A1 => n30741, A2 => n25891, B1 => n31089, B2 => 
                           n30734, ZN => n6777);
   U24646 : OAI22_X1 port map( A1 => n30741, A2 => n25890, B1 => n31092, B2 => 
                           n30734, ZN => n6778);
   U24647 : OAI22_X1 port map( A1 => n30741, A2 => n25889, B1 => n31095, B2 => 
                           n30734, ZN => n6779);
   U24648 : OAI22_X1 port map( A1 => n30742, A2 => n25888, B1 => n31098, B2 => 
                           n30734, ZN => n6780);
   U24649 : OAI22_X1 port map( A1 => n30742, A2 => n25887, B1 => n31101, B2 => 
                           n30734, ZN => n6781);
   U24650 : OAI22_X1 port map( A1 => n30742, A2 => n25886, B1 => n31104, B2 => 
                           n30734, ZN => n6782);
   U24651 : OAI22_X1 port map( A1 => n30742, A2 => n25885, B1 => n31107, B2 => 
                           n30734, ZN => n6783);
   U24652 : OAI22_X1 port map( A1 => n30742, A2 => n25884, B1 => n31110, B2 => 
                           n30734, ZN => n6784);
   U24653 : OAI22_X1 port map( A1 => n30742, A2 => n25883, B1 => n31113, B2 => 
                           n30734, ZN => n6785);
   U24654 : OAI22_X1 port map( A1 => n30742, A2 => n25882, B1 => n31116, B2 => 
                           n30734, ZN => n6786);
   U24655 : OAI22_X1 port map( A1 => n30742, A2 => n25881, B1 => n31119, B2 => 
                           n30734, ZN => n6787);
   U24656 : OAI22_X1 port map( A1 => n30742, A2 => n25880, B1 => n31122, B2 => 
                           n30734, ZN => n6788);
   U24657 : OAI22_X1 port map( A1 => n9672, A2 => n30762, B1 => n30945, B2 => 
                           n30756, ZN => n6857);
   U24658 : OAI22_X1 port map( A1 => n9671, A2 => n30762, B1 => n30948, B2 => 
                           n30756, ZN => n6858);
   U24659 : OAI22_X1 port map( A1 => n9670, A2 => n30762, B1 => n30951, B2 => 
                           n30756, ZN => n6859);
   U24660 : OAI22_X1 port map( A1 => n9669, A2 => n30762, B1 => n30954, B2 => 
                           n30756, ZN => n6860);
   U24661 : OAI22_X1 port map( A1 => n9668, A2 => n30762, B1 => n30957, B2 => 
                           n30756, ZN => n6861);
   U24662 : OAI22_X1 port map( A1 => n9667, A2 => n30762, B1 => n30960, B2 => 
                           n30756, ZN => n6862);
   U24663 : OAI22_X1 port map( A1 => n9666, A2 => n30762, B1 => n30963, B2 => 
                           n30756, ZN => n6863);
   U24664 : OAI22_X1 port map( A1 => n9665, A2 => n30762, B1 => n30966, B2 => 
                           n30756, ZN => n6864);
   U24665 : OAI22_X1 port map( A1 => n9664, A2 => n30762, B1 => n30969, B2 => 
                           n30756, ZN => n6865);
   U24666 : OAI22_X1 port map( A1 => n9663, A2 => n30762, B1 => n30972, B2 => 
                           n30756, ZN => n6866);
   U24667 : OAI22_X1 port map( A1 => n9662, A2 => n30762, B1 => n30975, B2 => 
                           n30756, ZN => n6867);
   U24668 : OAI22_X1 port map( A1 => n9661, A2 => n30763, B1 => n30978, B2 => 
                           n30756, ZN => n6868);
   U24669 : OAI22_X1 port map( A1 => n9660, A2 => n30763, B1 => n30981, B2 => 
                           n30757, ZN => n6869);
   U24670 : OAI22_X1 port map( A1 => n9659, A2 => n30763, B1 => n30984, B2 => 
                           n30757, ZN => n6870);
   U24671 : OAI22_X1 port map( A1 => n9658, A2 => n30763, B1 => n30987, B2 => 
                           n30757, ZN => n6871);
   U24672 : OAI22_X1 port map( A1 => n9657, A2 => n30763, B1 => n30990, B2 => 
                           n30757, ZN => n6872);
   U24673 : OAI22_X1 port map( A1 => n9656, A2 => n30763, B1 => n30993, B2 => 
                           n30757, ZN => n6873);
   U24674 : OAI22_X1 port map( A1 => n9655, A2 => n30763, B1 => n30996, B2 => 
                           n30757, ZN => n6874);
   U24675 : OAI22_X1 port map( A1 => n9654, A2 => n30763, B1 => n30999, B2 => 
                           n30757, ZN => n6875);
   U24676 : OAI22_X1 port map( A1 => n9653, A2 => n30763, B1 => n31002, B2 => 
                           n30757, ZN => n6876);
   U24677 : OAI22_X1 port map( A1 => n9652, A2 => n30763, B1 => n31005, B2 => 
                           n30757, ZN => n6877);
   U24678 : OAI22_X1 port map( A1 => n9651, A2 => n30763, B1 => n31008, B2 => 
                           n30757, ZN => n6878);
   U24679 : OAI22_X1 port map( A1 => n9650, A2 => n30763, B1 => n31011, B2 => 
                           n30757, ZN => n6879);
   U24680 : OAI22_X1 port map( A1 => n9649, A2 => n30764, B1 => n31014, B2 => 
                           n30757, ZN => n6880);
   U24681 : OAI22_X1 port map( A1 => n9648, A2 => n30764, B1 => n31017, B2 => 
                           n30758, ZN => n6881);
   U24682 : OAI22_X1 port map( A1 => n9647, A2 => n30764, B1 => n31020, B2 => 
                           n30758, ZN => n6882);
   U24683 : OAI22_X1 port map( A1 => n9646, A2 => n30764, B1 => n31023, B2 => 
                           n30758, ZN => n6883);
   U24684 : OAI22_X1 port map( A1 => n9645, A2 => n30764, B1 => n31026, B2 => 
                           n30758, ZN => n6884);
   U24685 : OAI22_X1 port map( A1 => n9644, A2 => n30764, B1 => n31029, B2 => 
                           n30758, ZN => n6885);
   U24686 : OAI22_X1 port map( A1 => n9643, A2 => n30764, B1 => n31032, B2 => 
                           n30758, ZN => n6886);
   U24687 : OAI22_X1 port map( A1 => n9642, A2 => n30764, B1 => n31035, B2 => 
                           n30758, ZN => n6887);
   U24688 : OAI22_X1 port map( A1 => n9641, A2 => n30764, B1 => n31038, B2 => 
                           n30758, ZN => n6888);
   U24689 : OAI22_X1 port map( A1 => n9640, A2 => n30764, B1 => n31041, B2 => 
                           n30758, ZN => n6889);
   U24690 : OAI22_X1 port map( A1 => n9639, A2 => n30764, B1 => n31044, B2 => 
                           n30758, ZN => n6890);
   U24691 : OAI22_X1 port map( A1 => n9638, A2 => n30764, B1 => n31047, B2 => 
                           n30758, ZN => n6891);
   U24692 : OAI22_X1 port map( A1 => n9637, A2 => n30765, B1 => n31050, B2 => 
                           n30758, ZN => n6892);
   U24693 : OAI22_X1 port map( A1 => n9636, A2 => n30765, B1 => n31053, B2 => 
                           n30759, ZN => n6893);
   U24694 : OAI22_X1 port map( A1 => n9635, A2 => n30765, B1 => n31056, B2 => 
                           n30759, ZN => n6894);
   U24695 : OAI22_X1 port map( A1 => n9634, A2 => n30765, B1 => n31059, B2 => 
                           n30759, ZN => n6895);
   U24696 : OAI22_X1 port map( A1 => n9633, A2 => n30765, B1 => n31062, B2 => 
                           n30759, ZN => n6896);
   U24697 : OAI22_X1 port map( A1 => n9632, A2 => n30765, B1 => n31065, B2 => 
                           n30759, ZN => n6897);
   U24698 : OAI22_X1 port map( A1 => n9631, A2 => n30765, B1 => n31068, B2 => 
                           n30759, ZN => n6898);
   U24699 : OAI22_X1 port map( A1 => n9630, A2 => n30765, B1 => n31071, B2 => 
                           n30759, ZN => n6899);
   U24700 : OAI22_X1 port map( A1 => n9629, A2 => n30765, B1 => n31074, B2 => 
                           n30759, ZN => n6900);
   U24701 : OAI22_X1 port map( A1 => n9628, A2 => n30765, B1 => n31077, B2 => 
                           n30759, ZN => n6901);
   U24702 : OAI22_X1 port map( A1 => n9627, A2 => n30765, B1 => n31080, B2 => 
                           n30759, ZN => n6902);
   U24703 : OAI22_X1 port map( A1 => n9626, A2 => n30765, B1 => n31083, B2 => 
                           n30759, ZN => n6903);
   U24704 : OAI22_X1 port map( A1 => n9625, A2 => n30766, B1 => n31086, B2 => 
                           n30759, ZN => n6904);
   U24705 : OAI22_X1 port map( A1 => n9624, A2 => n30766, B1 => n31089, B2 => 
                           n30760, ZN => n6905);
   U24706 : OAI22_X1 port map( A1 => n9623, A2 => n30766, B1 => n31092, B2 => 
                           n30760, ZN => n6906);
   U24707 : OAI22_X1 port map( A1 => n9622, A2 => n30766, B1 => n31095, B2 => 
                           n30760, ZN => n6907);
   U24708 : OAI22_X1 port map( A1 => n9621, A2 => n30766, B1 => n31098, B2 => 
                           n30760, ZN => n6908);
   U24709 : OAI22_X1 port map( A1 => n9620, A2 => n30766, B1 => n31101, B2 => 
                           n30760, ZN => n6909);
   U24710 : OAI22_X1 port map( A1 => n9619, A2 => n30766, B1 => n31104, B2 => 
                           n30760, ZN => n6910);
   U24711 : OAI22_X1 port map( A1 => n9618, A2 => n30766, B1 => n31107, B2 => 
                           n30760, ZN => n6911);
   U24712 : OAI22_X1 port map( A1 => n9617, A2 => n30766, B1 => n31110, B2 => 
                           n30760, ZN => n6912);
   U24713 : OAI22_X1 port map( A1 => n9616, A2 => n30766, B1 => n31113, B2 => 
                           n30760, ZN => n6913);
   U24714 : OAI22_X1 port map( A1 => n9615, A2 => n30766, B1 => n31116, B2 => 
                           n30760, ZN => n6914);
   U24715 : OAI22_X1 port map( A1 => n9614, A2 => n30766, B1 => n31119, B2 => 
                           n30760, ZN => n6915);
   U24716 : OAI22_X1 port map( A1 => n9613, A2 => n30767, B1 => n31122, B2 => 
                           n30760, ZN => n6916);
   U24717 : OAI22_X1 port map( A1 => n9286, A2 => n30812, B1 => n30945, B2 => 
                           n30806, ZN => n7113);
   U24718 : OAI22_X1 port map( A1 => n9281, A2 => n30812, B1 => n30948, B2 => 
                           n30806, ZN => n7114);
   U24719 : OAI22_X1 port map( A1 => n9276, A2 => n30812, B1 => n30951, B2 => 
                           n30806, ZN => n7115);
   U24720 : OAI22_X1 port map( A1 => n9271, A2 => n30812, B1 => n30954, B2 => 
                           n30806, ZN => n7116);
   U24721 : OAI22_X1 port map( A1 => n9266, A2 => n30812, B1 => n30957, B2 => 
                           n30806, ZN => n7117);
   U24722 : OAI22_X1 port map( A1 => n9261, A2 => n30812, B1 => n30960, B2 => 
                           n30806, ZN => n7118);
   U24723 : OAI22_X1 port map( A1 => n9256, A2 => n30812, B1 => n30963, B2 => 
                           n30806, ZN => n7119);
   U24724 : OAI22_X1 port map( A1 => n9251, A2 => n30812, B1 => n30966, B2 => 
                           n30806, ZN => n7120);
   U24725 : OAI22_X1 port map( A1 => n9246, A2 => n30812, B1 => n30969, B2 => 
                           n30806, ZN => n7121);
   U24726 : OAI22_X1 port map( A1 => n9241, A2 => n30812, B1 => n30972, B2 => 
                           n30806, ZN => n7122);
   U24727 : OAI22_X1 port map( A1 => n9236, A2 => n30812, B1 => n30975, B2 => 
                           n30806, ZN => n7123);
   U24728 : OAI22_X1 port map( A1 => n9231, A2 => n30813, B1 => n30978, B2 => 
                           n30806, ZN => n7124);
   U24729 : OAI22_X1 port map( A1 => n9226, A2 => n30813, B1 => n30981, B2 => 
                           n30807, ZN => n7125);
   U24730 : OAI22_X1 port map( A1 => n9221, A2 => n30813, B1 => n30984, B2 => 
                           n30807, ZN => n7126);
   U24731 : OAI22_X1 port map( A1 => n9216, A2 => n30813, B1 => n30987, B2 => 
                           n30807, ZN => n7127);
   U24732 : OAI22_X1 port map( A1 => n9211, A2 => n30813, B1 => n30990, B2 => 
                           n30807, ZN => n7128);
   U24733 : OAI22_X1 port map( A1 => n9206, A2 => n30813, B1 => n30993, B2 => 
                           n30807, ZN => n7129);
   U24734 : OAI22_X1 port map( A1 => n9201, A2 => n30813, B1 => n30996, B2 => 
                           n30807, ZN => n7130);
   U24735 : OAI22_X1 port map( A1 => n9196, A2 => n30813, B1 => n30999, B2 => 
                           n30807, ZN => n7131);
   U24736 : OAI22_X1 port map( A1 => n9191, A2 => n30813, B1 => n31002, B2 => 
                           n30807, ZN => n7132);
   U24737 : OAI22_X1 port map( A1 => n9186, A2 => n30813, B1 => n31005, B2 => 
                           n30807, ZN => n7133);
   U24738 : OAI22_X1 port map( A1 => n9181, A2 => n30813, B1 => n31008, B2 => 
                           n30807, ZN => n7134);
   U24739 : OAI22_X1 port map( A1 => n9176, A2 => n30813, B1 => n31011, B2 => 
                           n30807, ZN => n7135);
   U24740 : OAI22_X1 port map( A1 => n9171, A2 => n30814, B1 => n31014, B2 => 
                           n30807, ZN => n7136);
   U24741 : OAI22_X1 port map( A1 => n9166, A2 => n30814, B1 => n31017, B2 => 
                           n30808, ZN => n7137);
   U24742 : OAI22_X1 port map( A1 => n9161, A2 => n30814, B1 => n31020, B2 => 
                           n30808, ZN => n7138);
   U24743 : OAI22_X1 port map( A1 => n9156, A2 => n30814, B1 => n31023, B2 => 
                           n30808, ZN => n7139);
   U24744 : OAI22_X1 port map( A1 => n9151, A2 => n30814, B1 => n31026, B2 => 
                           n30808, ZN => n7140);
   U24745 : OAI22_X1 port map( A1 => n9146, A2 => n30814, B1 => n31029, B2 => 
                           n30808, ZN => n7141);
   U24746 : OAI22_X1 port map( A1 => n9141, A2 => n30814, B1 => n31032, B2 => 
                           n30808, ZN => n7142);
   U24747 : OAI22_X1 port map( A1 => n9136, A2 => n30814, B1 => n31035, B2 => 
                           n30808, ZN => n7143);
   U24748 : OAI22_X1 port map( A1 => n9131, A2 => n30814, B1 => n31038, B2 => 
                           n30808, ZN => n7144);
   U24749 : OAI22_X1 port map( A1 => n9126, A2 => n30814, B1 => n31041, B2 => 
                           n30808, ZN => n7145);
   U24750 : OAI22_X1 port map( A1 => n9121, A2 => n30814, B1 => n31044, B2 => 
                           n30808, ZN => n7146);
   U24751 : OAI22_X1 port map( A1 => n9116, A2 => n30814, B1 => n31047, B2 => 
                           n30808, ZN => n7147);
   U24752 : OAI22_X1 port map( A1 => n9111, A2 => n30815, B1 => n31050, B2 => 
                           n30808, ZN => n7148);
   U24753 : OAI22_X1 port map( A1 => n9106, A2 => n30815, B1 => n31053, B2 => 
                           n30809, ZN => n7149);
   U24754 : OAI22_X1 port map( A1 => n9101, A2 => n30815, B1 => n31056, B2 => 
                           n30809, ZN => n7150);
   U24755 : OAI22_X1 port map( A1 => n9096, A2 => n30815, B1 => n31059, B2 => 
                           n30809, ZN => n7151);
   U24756 : OAI22_X1 port map( A1 => n9091, A2 => n30815, B1 => n31062, B2 => 
                           n30809, ZN => n7152);
   U24757 : OAI22_X1 port map( A1 => n9086, A2 => n30815, B1 => n31065, B2 => 
                           n30809, ZN => n7153);
   U24758 : OAI22_X1 port map( A1 => n9081, A2 => n30815, B1 => n31068, B2 => 
                           n30809, ZN => n7154);
   U24759 : OAI22_X1 port map( A1 => n9076, A2 => n30815, B1 => n31071, B2 => 
                           n30809, ZN => n7155);
   U24760 : OAI22_X1 port map( A1 => n9071, A2 => n30815, B1 => n31074, B2 => 
                           n30809, ZN => n7156);
   U24761 : OAI22_X1 port map( A1 => n9066, A2 => n30815, B1 => n31077, B2 => 
                           n30809, ZN => n7157);
   U24762 : OAI22_X1 port map( A1 => n9061, A2 => n30815, B1 => n31080, B2 => 
                           n30809, ZN => n7158);
   U24763 : OAI22_X1 port map( A1 => n9056, A2 => n30815, B1 => n31083, B2 => 
                           n30809, ZN => n7159);
   U24764 : OAI22_X1 port map( A1 => n9051, A2 => n30816, B1 => n31086, B2 => 
                           n30809, ZN => n7160);
   U24765 : OAI22_X1 port map( A1 => n9046, A2 => n30816, B1 => n31089, B2 => 
                           n30810, ZN => n7161);
   U24766 : OAI22_X1 port map( A1 => n9041, A2 => n30816, B1 => n31092, B2 => 
                           n30810, ZN => n7162);
   U24767 : OAI22_X1 port map( A1 => n9036, A2 => n30816, B1 => n31095, B2 => 
                           n30810, ZN => n7163);
   U24768 : OAI22_X1 port map( A1 => n9031, A2 => n30816, B1 => n31098, B2 => 
                           n30810, ZN => n7164);
   U24769 : OAI22_X1 port map( A1 => n9026, A2 => n30816, B1 => n31101, B2 => 
                           n30810, ZN => n7165);
   U24770 : OAI22_X1 port map( A1 => n9021, A2 => n30816, B1 => n31104, B2 => 
                           n30810, ZN => n7166);
   U24771 : OAI22_X1 port map( A1 => n9016, A2 => n30816, B1 => n31107, B2 => 
                           n30810, ZN => n7167);
   U24772 : OAI22_X1 port map( A1 => n9011, A2 => n30816, B1 => n31110, B2 => 
                           n30810, ZN => n7168);
   U24773 : OAI22_X1 port map( A1 => n9006, A2 => n30816, B1 => n31113, B2 => 
                           n30810, ZN => n7169);
   U24774 : OAI22_X1 port map( A1 => n9001, A2 => n30816, B1 => n31116, B2 => 
                           n30810, ZN => n7170);
   U24775 : OAI22_X1 port map( A1 => n8996, A2 => n30816, B1 => n31119, B2 => 
                           n30810, ZN => n7171);
   U24776 : OAI22_X1 port map( A1 => n8991, A2 => n30817, B1 => n31122, B2 => 
                           n30810, ZN => n7172);
   U24777 : OAI22_X1 port map( A1 => n9999, A2 => n30828, B1 => n30977, B2 => 
                           n30818, ZN => n7188);
   U24778 : OAI22_X1 port map( A1 => n9994, A2 => n30828, B1 => n30980, B2 => 
                           n30819, ZN => n7189);
   U24779 : OAI22_X1 port map( A1 => n9989, A2 => n30828, B1 => n30983, B2 => 
                           n30819, ZN => n7190);
   U24780 : OAI22_X1 port map( A1 => n9984, A2 => n30828, B1 => n30986, B2 => 
                           n30819, ZN => n7191);
   U24781 : OAI22_X1 port map( A1 => n9979, A2 => n30828, B1 => n30989, B2 => 
                           n30819, ZN => n7192);
   U24782 : OAI22_X1 port map( A1 => n9974, A2 => n30828, B1 => n30992, B2 => 
                           n30819, ZN => n7193);
   U24783 : OAI22_X1 port map( A1 => n9969, A2 => n30827, B1 => n30995, B2 => 
                           n30819, ZN => n7194);
   U24784 : OAI22_X1 port map( A1 => n9964, A2 => n30827, B1 => n30998, B2 => 
                           n30819, ZN => n7195);
   U24785 : OAI22_X1 port map( A1 => n9959, A2 => n30827, B1 => n31001, B2 => 
                           n30819, ZN => n7196);
   U24786 : OAI22_X1 port map( A1 => n9954, A2 => n30827, B1 => n31004, B2 => 
                           n30819, ZN => n7197);
   U24787 : OAI22_X1 port map( A1 => n9949, A2 => n30827, B1 => n31007, B2 => 
                           n30819, ZN => n7198);
   U24788 : OAI22_X1 port map( A1 => n9944, A2 => n30827, B1 => n31010, B2 => 
                           n30819, ZN => n7199);
   U24789 : OAI22_X1 port map( A1 => n9939, A2 => n30827, B1 => n31013, B2 => 
                           n30819, ZN => n7200);
   U24790 : OAI22_X1 port map( A1 => n9934, A2 => n30827, B1 => n31016, B2 => 
                           n30820, ZN => n7201);
   U24791 : OAI22_X1 port map( A1 => n9929, A2 => n30827, B1 => n31019, B2 => 
                           n30820, ZN => n7202);
   U24792 : OAI22_X1 port map( A1 => n9924, A2 => n30827, B1 => n31022, B2 => 
                           n30820, ZN => n7203);
   U24793 : OAI22_X1 port map( A1 => n9919, A2 => n30827, B1 => n31025, B2 => 
                           n30820, ZN => n7204);
   U24794 : OAI22_X1 port map( A1 => n9914, A2 => n30827, B1 => n31028, B2 => 
                           n30820, ZN => n7205);
   U24795 : OAI22_X1 port map( A1 => n9909, A2 => n30826, B1 => n31031, B2 => 
                           n30820, ZN => n7206);
   U24796 : OAI22_X1 port map( A1 => n9904, A2 => n30826, B1 => n31034, B2 => 
                           n30820, ZN => n7207);
   U24797 : OAI22_X1 port map( A1 => n9899, A2 => n30826, B1 => n31037, B2 => 
                           n30820, ZN => n7208);
   U24798 : OAI22_X1 port map( A1 => n9894, A2 => n30826, B1 => n31040, B2 => 
                           n30820, ZN => n7209);
   U24799 : OAI22_X1 port map( A1 => n9889, A2 => n30826, B1 => n31043, B2 => 
                           n30820, ZN => n7210);
   U24800 : OAI22_X1 port map( A1 => n9884, A2 => n30826, B1 => n31046, B2 => 
                           n30820, ZN => n7211);
   U24801 : OAI22_X1 port map( A1 => n9879, A2 => n30826, B1 => n31049, B2 => 
                           n30820, ZN => n7212);
   U24802 : OAI22_X1 port map( A1 => n9874, A2 => n30826, B1 => n31052, B2 => 
                           n30821, ZN => n7213);
   U24803 : OAI22_X1 port map( A1 => n9869, A2 => n30826, B1 => n31055, B2 => 
                           n30821, ZN => n7214);
   U24804 : OAI22_X1 port map( A1 => n9864, A2 => n30826, B1 => n31058, B2 => 
                           n30821, ZN => n7215);
   U24805 : OAI22_X1 port map( A1 => n9859, A2 => n30826, B1 => n31061, B2 => 
                           n30821, ZN => n7216);
   U24806 : OAI22_X1 port map( A1 => n9854, A2 => n30825, B1 => n31064, B2 => 
                           n30821, ZN => n7217);
   U24807 : OAI22_X1 port map( A1 => n9849, A2 => n30825, B1 => n31067, B2 => 
                           n30821, ZN => n7218);
   U24808 : OAI22_X1 port map( A1 => n9844, A2 => n30825, B1 => n31070, B2 => 
                           n30821, ZN => n7219);
   U24809 : OAI22_X1 port map( A1 => n9839, A2 => n30825, B1 => n31073, B2 => 
                           n30821, ZN => n7220);
   U24810 : OAI22_X1 port map( A1 => n9834, A2 => n30825, B1 => n31076, B2 => 
                           n30821, ZN => n7221);
   U24811 : OAI22_X1 port map( A1 => n9829, A2 => n30825, B1 => n31079, B2 => 
                           n30821, ZN => n7222);
   U24812 : OAI22_X1 port map( A1 => n9824, A2 => n30825, B1 => n31082, B2 => 
                           n30821, ZN => n7223);
   U24813 : OAI22_X1 port map( A1 => n9819, A2 => n30825, B1 => n31085, B2 => 
                           n30821, ZN => n7224);
   U24814 : OAI22_X1 port map( A1 => n9814, A2 => n30825, B1 => n31088, B2 => 
                           n30822, ZN => n7225);
   U24815 : OAI22_X1 port map( A1 => n9809, A2 => n30825, B1 => n31091, B2 => 
                           n30822, ZN => n7226);
   U24816 : OAI22_X1 port map( A1 => n9804, A2 => n30825, B1 => n31094, B2 => 
                           n30822, ZN => n7227);
   U24817 : OAI22_X1 port map( A1 => n9799, A2 => n30825, B1 => n31097, B2 => 
                           n30822, ZN => n7228);
   U24818 : OAI22_X1 port map( A1 => n9794, A2 => n30824, B1 => n31100, B2 => 
                           n30822, ZN => n7229);
   U24819 : OAI22_X1 port map( A1 => n9789, A2 => n30824, B1 => n31103, B2 => 
                           n30822, ZN => n7230);
   U24820 : OAI22_X1 port map( A1 => n9784, A2 => n30824, B1 => n31106, B2 => 
                           n30822, ZN => n7231);
   U24821 : OAI22_X1 port map( A1 => n9779, A2 => n30824, B1 => n31109, B2 => 
                           n30822, ZN => n7232);
   U24822 : OAI22_X1 port map( A1 => n9774, A2 => n30824, B1 => n31112, B2 => 
                           n30822, ZN => n7233);
   U24823 : OAI22_X1 port map( A1 => n9769, A2 => n30824, B1 => n31115, B2 => 
                           n30822, ZN => n7234);
   U24824 : OAI22_X1 port map( A1 => n9764, A2 => n30824, B1 => n31118, B2 => 
                           n30822, ZN => n7235);
   U24825 : OAI22_X1 port map( A1 => n9759, A2 => n30824, B1 => n31121, B2 => 
                           n30822, ZN => n7236);
   U24826 : OAI22_X1 port map( A1 => n30838, A2 => n25653, B1 => n30944, B2 => 
                           n30830, ZN => n7241);
   U24827 : OAI22_X1 port map( A1 => n30838, A2 => n25652, B1 => n30947, B2 => 
                           n30830, ZN => n7242);
   U24828 : OAI22_X1 port map( A1 => n30838, A2 => n25651, B1 => n30950, B2 => 
                           n30830, ZN => n7243);
   U24829 : OAI22_X1 port map( A1 => n30838, A2 => n25650, B1 => n30953, B2 => 
                           n30830, ZN => n7244);
   U24830 : OAI22_X1 port map( A1 => n30838, A2 => n25649, B1 => n30956, B2 => 
                           n30830, ZN => n7245);
   U24831 : OAI22_X1 port map( A1 => n30838, A2 => n25648, B1 => n30959, B2 => 
                           n30830, ZN => n7246);
   U24832 : OAI22_X1 port map( A1 => n30838, A2 => n25647, B1 => n30962, B2 => 
                           n30830, ZN => n7247);
   U24833 : OAI22_X1 port map( A1 => n30838, A2 => n25646, B1 => n30965, B2 => 
                           n30830, ZN => n7248);
   U24834 : OAI22_X1 port map( A1 => n30838, A2 => n25645, B1 => n30968, B2 => 
                           n30830, ZN => n7249);
   U24835 : OAI22_X1 port map( A1 => n30838, A2 => n25644, B1 => n30971, B2 => 
                           n30830, ZN => n7250);
   U24836 : OAI22_X1 port map( A1 => n30838, A2 => n25643, B1 => n30974, B2 => 
                           n30830, ZN => n7251);
   U24837 : OAI22_X1 port map( A1 => n30838, A2 => n25642, B1 => n30977, B2 => 
                           n30830, ZN => n7252);
   U24838 : OAI22_X1 port map( A1 => n30839, A2 => n25641, B1 => n30980, B2 => 
                           n30831, ZN => n7253);
   U24839 : OAI22_X1 port map( A1 => n30839, A2 => n25640, B1 => n30983, B2 => 
                           n30831, ZN => n7254);
   U24840 : OAI22_X1 port map( A1 => n30839, A2 => n25639, B1 => n30986, B2 => 
                           n30831, ZN => n7255);
   U24841 : OAI22_X1 port map( A1 => n30839, A2 => n25638, B1 => n30989, B2 => 
                           n30831, ZN => n7256);
   U24842 : OAI22_X1 port map( A1 => n30839, A2 => n25637, B1 => n30992, B2 => 
                           n30831, ZN => n7257);
   U24843 : OAI22_X1 port map( A1 => n30839, A2 => n25636, B1 => n30995, B2 => 
                           n30831, ZN => n7258);
   U24844 : OAI22_X1 port map( A1 => n30839, A2 => n25635, B1 => n30998, B2 => 
                           n30831, ZN => n7259);
   U24845 : OAI22_X1 port map( A1 => n30839, A2 => n25634, B1 => n31001, B2 => 
                           n30831, ZN => n7260);
   U24846 : OAI22_X1 port map( A1 => n30839, A2 => n25633, B1 => n31004, B2 => 
                           n30831, ZN => n7261);
   U24847 : OAI22_X1 port map( A1 => n30839, A2 => n25632, B1 => n31007, B2 => 
                           n30831, ZN => n7262);
   U24848 : OAI22_X1 port map( A1 => n30839, A2 => n25631, B1 => n31010, B2 => 
                           n30831, ZN => n7263);
   U24849 : OAI22_X1 port map( A1 => n30839, A2 => n25630, B1 => n31013, B2 => 
                           n30831, ZN => n7264);
   U24850 : OAI22_X1 port map( A1 => n30839, A2 => n25629, B1 => n31016, B2 => 
                           n30832, ZN => n7265);
   U24851 : OAI22_X1 port map( A1 => n30840, A2 => n25628, B1 => n31019, B2 => 
                           n30832, ZN => n7266);
   U24852 : OAI22_X1 port map( A1 => n30840, A2 => n25627, B1 => n31022, B2 => 
                           n30832, ZN => n7267);
   U24853 : OAI22_X1 port map( A1 => n30840, A2 => n25626, B1 => n31025, B2 => 
                           n30832, ZN => n7268);
   U24854 : OAI22_X1 port map( A1 => n30840, A2 => n25625, B1 => n31028, B2 => 
                           n30832, ZN => n7269);
   U24855 : OAI22_X1 port map( A1 => n30840, A2 => n25624, B1 => n31031, B2 => 
                           n30832, ZN => n7270);
   U24856 : OAI22_X1 port map( A1 => n30840, A2 => n25623, B1 => n31034, B2 => 
                           n30832, ZN => n7271);
   U24857 : OAI22_X1 port map( A1 => n30840, A2 => n25622, B1 => n31037, B2 => 
                           n30832, ZN => n7272);
   U24858 : OAI22_X1 port map( A1 => n30840, A2 => n25621, B1 => n31040, B2 => 
                           n30832, ZN => n7273);
   U24859 : OAI22_X1 port map( A1 => n30840, A2 => n25620, B1 => n31043, B2 => 
                           n30832, ZN => n7274);
   U24860 : OAI22_X1 port map( A1 => n30840, A2 => n25619, B1 => n31046, B2 => 
                           n30832, ZN => n7275);
   U24861 : OAI22_X1 port map( A1 => n30840, A2 => n25618, B1 => n31049, B2 => 
                           n30832, ZN => n7276);
   U24862 : OAI22_X1 port map( A1 => n30840, A2 => n25617, B1 => n31052, B2 => 
                           n30833, ZN => n7277);
   U24863 : OAI22_X1 port map( A1 => n30840, A2 => n25616, B1 => n31055, B2 => 
                           n30833, ZN => n7278);
   U24864 : OAI22_X1 port map( A1 => n30841, A2 => n25615, B1 => n31058, B2 => 
                           n30833, ZN => n7279);
   U24865 : OAI22_X1 port map( A1 => n30841, A2 => n25614, B1 => n31061, B2 => 
                           n30833, ZN => n7280);
   U24866 : OAI22_X1 port map( A1 => n30841, A2 => n25613, B1 => n31064, B2 => 
                           n30833, ZN => n7281);
   U24867 : OAI22_X1 port map( A1 => n30841, A2 => n25612, B1 => n31067, B2 => 
                           n30833, ZN => n7282);
   U24868 : OAI22_X1 port map( A1 => n30841, A2 => n25611, B1 => n31070, B2 => 
                           n30833, ZN => n7283);
   U24869 : OAI22_X1 port map( A1 => n30841, A2 => n25610, B1 => n31073, B2 => 
                           n30833, ZN => n7284);
   U24870 : OAI22_X1 port map( A1 => n30841, A2 => n25609, B1 => n31076, B2 => 
                           n30833, ZN => n7285);
   U24871 : OAI22_X1 port map( A1 => n30841, A2 => n25608, B1 => n31079, B2 => 
                           n30833, ZN => n7286);
   U24872 : OAI22_X1 port map( A1 => n30841, A2 => n25607, B1 => n31082, B2 => 
                           n30833, ZN => n7287);
   U24873 : OAI22_X1 port map( A1 => n30841, A2 => n25606, B1 => n31085, B2 => 
                           n30833, ZN => n7288);
   U24874 : OAI22_X1 port map( A1 => n30841, A2 => n25605, B1 => n31088, B2 => 
                           n30834, ZN => n7289);
   U24875 : OAI22_X1 port map( A1 => n30841, A2 => n25604, B1 => n31091, B2 => 
                           n30834, ZN => n7290);
   U24876 : OAI22_X1 port map( A1 => n30841, A2 => n25603, B1 => n31094, B2 => 
                           n30834, ZN => n7291);
   U24877 : OAI22_X1 port map( A1 => n30842, A2 => n25602, B1 => n31097, B2 => 
                           n30834, ZN => n7292);
   U24878 : OAI22_X1 port map( A1 => n30842, A2 => n25601, B1 => n31100, B2 => 
                           n30834, ZN => n7293);
   U24879 : OAI22_X1 port map( A1 => n30842, A2 => n25600, B1 => n31103, B2 => 
                           n30834, ZN => n7294);
   U24880 : OAI22_X1 port map( A1 => n30842, A2 => n25599, B1 => n31106, B2 => 
                           n30834, ZN => n7295);
   U24881 : OAI22_X1 port map( A1 => n30842, A2 => n25598, B1 => n31109, B2 => 
                           n30834, ZN => n7296);
   U24882 : OAI22_X1 port map( A1 => n30842, A2 => n25597, B1 => n31112, B2 => 
                           n30834, ZN => n7297);
   U24883 : OAI22_X1 port map( A1 => n30842, A2 => n25596, B1 => n31115, B2 => 
                           n30834, ZN => n7298);
   U24884 : OAI22_X1 port map( A1 => n30842, A2 => n25595, B1 => n31118, B2 => 
                           n30834, ZN => n7299);
   U24885 : OAI22_X1 port map( A1 => n30842, A2 => n25594, B1 => n31121, B2 => 
                           n30834, ZN => n7300);
   U24886 : OAI22_X1 port map( A1 => n30864, A2 => n25520, B1 => n30944, B2 => 
                           n30856, ZN => n7369);
   U24887 : OAI22_X1 port map( A1 => n30864, A2 => n25519, B1 => n30947, B2 => 
                           n30856, ZN => n7370);
   U24888 : OAI22_X1 port map( A1 => n30864, A2 => n25518, B1 => n30950, B2 => 
                           n30856, ZN => n7371);
   U24889 : OAI22_X1 port map( A1 => n30864, A2 => n25517, B1 => n30953, B2 => 
                           n30856, ZN => n7372);
   U24890 : OAI22_X1 port map( A1 => n30864, A2 => n25516, B1 => n30956, B2 => 
                           n30856, ZN => n7373);
   U24891 : OAI22_X1 port map( A1 => n30864, A2 => n25515, B1 => n30959, B2 => 
                           n30856, ZN => n7374);
   U24892 : OAI22_X1 port map( A1 => n30864, A2 => n25514, B1 => n30962, B2 => 
                           n30856, ZN => n7375);
   U24893 : OAI22_X1 port map( A1 => n30864, A2 => n25513, B1 => n30965, B2 => 
                           n30856, ZN => n7376);
   U24894 : OAI22_X1 port map( A1 => n30864, A2 => n25512, B1 => n30968, B2 => 
                           n30856, ZN => n7377);
   U24895 : OAI22_X1 port map( A1 => n30864, A2 => n25511, B1 => n30971, B2 => 
                           n30856, ZN => n7378);
   U24896 : OAI22_X1 port map( A1 => n30864, A2 => n25510, B1 => n30974, B2 => 
                           n30856, ZN => n7379);
   U24897 : OAI22_X1 port map( A1 => n30864, A2 => n25509, B1 => n30977, B2 => 
                           n30856, ZN => n7380);
   U24898 : OAI22_X1 port map( A1 => n30865, A2 => n25508, B1 => n30980, B2 => 
                           n30857, ZN => n7381);
   U24899 : OAI22_X1 port map( A1 => n30865, A2 => n25507, B1 => n30983, B2 => 
                           n30857, ZN => n7382);
   U24900 : OAI22_X1 port map( A1 => n30865, A2 => n25506, B1 => n30986, B2 => 
                           n30857, ZN => n7383);
   U24901 : OAI22_X1 port map( A1 => n30865, A2 => n25505, B1 => n30989, B2 => 
                           n30857, ZN => n7384);
   U24902 : OAI22_X1 port map( A1 => n30865, A2 => n25504, B1 => n30992, B2 => 
                           n30857, ZN => n7385);
   U24903 : OAI22_X1 port map( A1 => n30865, A2 => n25503, B1 => n30995, B2 => 
                           n30857, ZN => n7386);
   U24904 : OAI22_X1 port map( A1 => n30865, A2 => n25502, B1 => n30998, B2 => 
                           n30857, ZN => n7387);
   U24905 : OAI22_X1 port map( A1 => n30865, A2 => n25501, B1 => n31001, B2 => 
                           n30857, ZN => n7388);
   U24906 : OAI22_X1 port map( A1 => n30865, A2 => n25500, B1 => n31004, B2 => 
                           n30857, ZN => n7389);
   U24907 : OAI22_X1 port map( A1 => n30865, A2 => n25499, B1 => n31007, B2 => 
                           n30857, ZN => n7390);
   U24908 : OAI22_X1 port map( A1 => n30865, A2 => n25498, B1 => n31010, B2 => 
                           n30857, ZN => n7391);
   U24909 : OAI22_X1 port map( A1 => n30865, A2 => n25497, B1 => n31013, B2 => 
                           n30857, ZN => n7392);
   U24910 : OAI22_X1 port map( A1 => n30865, A2 => n25496, B1 => n31016, B2 => 
                           n30858, ZN => n7393);
   U24911 : OAI22_X1 port map( A1 => n30866, A2 => n25495, B1 => n31019, B2 => 
                           n30858, ZN => n7394);
   U24912 : OAI22_X1 port map( A1 => n30866, A2 => n25494, B1 => n31022, B2 => 
                           n30858, ZN => n7395);
   U24913 : OAI22_X1 port map( A1 => n30866, A2 => n25493, B1 => n31025, B2 => 
                           n30858, ZN => n7396);
   U24914 : OAI22_X1 port map( A1 => n30866, A2 => n25492, B1 => n31028, B2 => 
                           n30858, ZN => n7397);
   U24915 : OAI22_X1 port map( A1 => n30866, A2 => n25491, B1 => n31031, B2 => 
                           n30858, ZN => n7398);
   U24916 : OAI22_X1 port map( A1 => n30866, A2 => n25490, B1 => n31034, B2 => 
                           n30858, ZN => n7399);
   U24917 : OAI22_X1 port map( A1 => n30866, A2 => n25489, B1 => n31037, B2 => 
                           n30858, ZN => n7400);
   U24918 : OAI22_X1 port map( A1 => n30866, A2 => n25488, B1 => n31040, B2 => 
                           n30858, ZN => n7401);
   U24919 : OAI22_X1 port map( A1 => n30866, A2 => n25487, B1 => n31043, B2 => 
                           n30858, ZN => n7402);
   U24920 : OAI22_X1 port map( A1 => n30866, A2 => n25486, B1 => n31046, B2 => 
                           n30858, ZN => n7403);
   U24921 : OAI22_X1 port map( A1 => n30866, A2 => n25485, B1 => n31049, B2 => 
                           n30858, ZN => n7404);
   U24922 : OAI22_X1 port map( A1 => n30866, A2 => n25484, B1 => n31052, B2 => 
                           n30859, ZN => n7405);
   U24923 : OAI22_X1 port map( A1 => n30866, A2 => n25483, B1 => n31055, B2 => 
                           n30859, ZN => n7406);
   U24924 : OAI22_X1 port map( A1 => n30867, A2 => n25482, B1 => n31058, B2 => 
                           n30859, ZN => n7407);
   U24925 : OAI22_X1 port map( A1 => n30867, A2 => n25481, B1 => n31061, B2 => 
                           n30859, ZN => n7408);
   U24926 : OAI22_X1 port map( A1 => n30867, A2 => n25480, B1 => n31064, B2 => 
                           n30859, ZN => n7409);
   U24927 : OAI22_X1 port map( A1 => n30867, A2 => n25479, B1 => n31067, B2 => 
                           n30859, ZN => n7410);
   U24928 : OAI22_X1 port map( A1 => n30867, A2 => n25478, B1 => n31070, B2 => 
                           n30859, ZN => n7411);
   U24929 : OAI22_X1 port map( A1 => n30867, A2 => n25477, B1 => n31073, B2 => 
                           n30859, ZN => n7412);
   U24930 : OAI22_X1 port map( A1 => n30867, A2 => n25476, B1 => n31076, B2 => 
                           n30859, ZN => n7413);
   U24931 : OAI22_X1 port map( A1 => n30867, A2 => n25475, B1 => n31079, B2 => 
                           n30859, ZN => n7414);
   U24932 : OAI22_X1 port map( A1 => n30867, A2 => n25474, B1 => n31082, B2 => 
                           n30859, ZN => n7415);
   U24933 : OAI22_X1 port map( A1 => n30867, A2 => n25473, B1 => n31085, B2 => 
                           n30859, ZN => n7416);
   U24934 : OAI22_X1 port map( A1 => n30867, A2 => n25472, B1 => n31088, B2 => 
                           n30860, ZN => n7417);
   U24935 : OAI22_X1 port map( A1 => n30867, A2 => n25471, B1 => n31091, B2 => 
                           n30860, ZN => n7418);
   U24936 : OAI22_X1 port map( A1 => n30867, A2 => n25470, B1 => n31094, B2 => 
                           n30860, ZN => n7419);
   U24937 : OAI22_X1 port map( A1 => n30868, A2 => n25469, B1 => n31097, B2 => 
                           n30860, ZN => n7420);
   U24938 : OAI22_X1 port map( A1 => n30868, A2 => n25468, B1 => n31100, B2 => 
                           n30860, ZN => n7421);
   U24939 : OAI22_X1 port map( A1 => n30868, A2 => n25467, B1 => n31103, B2 => 
                           n30860, ZN => n7422);
   U24940 : OAI22_X1 port map( A1 => n30868, A2 => n25466, B1 => n31106, B2 => 
                           n30860, ZN => n7423);
   U24941 : OAI22_X1 port map( A1 => n30868, A2 => n25465, B1 => n31109, B2 => 
                           n30860, ZN => n7424);
   U24942 : OAI22_X1 port map( A1 => n30868, A2 => n25464, B1 => n31112, B2 => 
                           n30860, ZN => n7425);
   U24943 : OAI22_X1 port map( A1 => n30868, A2 => n25463, B1 => n31115, B2 => 
                           n30860, ZN => n7426);
   U24944 : OAI22_X1 port map( A1 => n30868, A2 => n25462, B1 => n31118, B2 => 
                           n30860, ZN => n7427);
   U24945 : OAI22_X1 port map( A1 => n30868, A2 => n25461, B1 => n31121, B2 => 
                           n30860, ZN => n7428);
   U24946 : OAI22_X1 port map( A1 => n9285, A2 => n30888, B1 => n30944, B2 => 
                           n30882, ZN => n7497);
   U24947 : OAI22_X1 port map( A1 => n9280, A2 => n30888, B1 => n30947, B2 => 
                           n30882, ZN => n7498);
   U24948 : OAI22_X1 port map( A1 => n9275, A2 => n30888, B1 => n30950, B2 => 
                           n30882, ZN => n7499);
   U24949 : OAI22_X1 port map( A1 => n9270, A2 => n30888, B1 => n30953, B2 => 
                           n30882, ZN => n7500);
   U24950 : OAI22_X1 port map( A1 => n9265, A2 => n30888, B1 => n30956, B2 => 
                           n30882, ZN => n7501);
   U24951 : OAI22_X1 port map( A1 => n9260, A2 => n30888, B1 => n30959, B2 => 
                           n30882, ZN => n7502);
   U24952 : OAI22_X1 port map( A1 => n9255, A2 => n30888, B1 => n30962, B2 => 
                           n30882, ZN => n7503);
   U24953 : OAI22_X1 port map( A1 => n9250, A2 => n30888, B1 => n30965, B2 => 
                           n30882, ZN => n7504);
   U24954 : OAI22_X1 port map( A1 => n9245, A2 => n30888, B1 => n30968, B2 => 
                           n30882, ZN => n7505);
   U24955 : OAI22_X1 port map( A1 => n9240, A2 => n30888, B1 => n30971, B2 => 
                           n30882, ZN => n7506);
   U24956 : OAI22_X1 port map( A1 => n9235, A2 => n30888, B1 => n30974, B2 => 
                           n30882, ZN => n7507);
   U24957 : OAI22_X1 port map( A1 => n9230, A2 => n30889, B1 => n30977, B2 => 
                           n30882, ZN => n7508);
   U24958 : OAI22_X1 port map( A1 => n9225, A2 => n30889, B1 => n30980, B2 => 
                           n30883, ZN => n7509);
   U24959 : OAI22_X1 port map( A1 => n9220, A2 => n30889, B1 => n30983, B2 => 
                           n30883, ZN => n7510);
   U24960 : OAI22_X1 port map( A1 => n9215, A2 => n30889, B1 => n30986, B2 => 
                           n30883, ZN => n7511);
   U24961 : OAI22_X1 port map( A1 => n9210, A2 => n30889, B1 => n30989, B2 => 
                           n30883, ZN => n7512);
   U24962 : OAI22_X1 port map( A1 => n9205, A2 => n30889, B1 => n30992, B2 => 
                           n30883, ZN => n7513);
   U24963 : OAI22_X1 port map( A1 => n9200, A2 => n30889, B1 => n30995, B2 => 
                           n30883, ZN => n7514);
   U24964 : OAI22_X1 port map( A1 => n9195, A2 => n30889, B1 => n30998, B2 => 
                           n30883, ZN => n7515);
   U24965 : OAI22_X1 port map( A1 => n9190, A2 => n30889, B1 => n31001, B2 => 
                           n30883, ZN => n7516);
   U24966 : OAI22_X1 port map( A1 => n9185, A2 => n30889, B1 => n31004, B2 => 
                           n30883, ZN => n7517);
   U24967 : OAI22_X1 port map( A1 => n9180, A2 => n30889, B1 => n31007, B2 => 
                           n30883, ZN => n7518);
   U24968 : OAI22_X1 port map( A1 => n9175, A2 => n30889, B1 => n31010, B2 => 
                           n30883, ZN => n7519);
   U24969 : OAI22_X1 port map( A1 => n9170, A2 => n30890, B1 => n31013, B2 => 
                           n30883, ZN => n7520);
   U24970 : OAI22_X1 port map( A1 => n9165, A2 => n30890, B1 => n31016, B2 => 
                           n30884, ZN => n7521);
   U24971 : OAI22_X1 port map( A1 => n9160, A2 => n30890, B1 => n31019, B2 => 
                           n30884, ZN => n7522);
   U24972 : OAI22_X1 port map( A1 => n9155, A2 => n30890, B1 => n31022, B2 => 
                           n30884, ZN => n7523);
   U24973 : OAI22_X1 port map( A1 => n9150, A2 => n30890, B1 => n31025, B2 => 
                           n30884, ZN => n7524);
   U24974 : OAI22_X1 port map( A1 => n9145, A2 => n30890, B1 => n31028, B2 => 
                           n30884, ZN => n7525);
   U24975 : OAI22_X1 port map( A1 => n9140, A2 => n30890, B1 => n31031, B2 => 
                           n30884, ZN => n7526);
   U24976 : OAI22_X1 port map( A1 => n9135, A2 => n30890, B1 => n31034, B2 => 
                           n30884, ZN => n7527);
   U24977 : OAI22_X1 port map( A1 => n9130, A2 => n30890, B1 => n31037, B2 => 
                           n30884, ZN => n7528);
   U24978 : OAI22_X1 port map( A1 => n9125, A2 => n30890, B1 => n31040, B2 => 
                           n30884, ZN => n7529);
   U24979 : OAI22_X1 port map( A1 => n9120, A2 => n30890, B1 => n31043, B2 => 
                           n30884, ZN => n7530);
   U24980 : OAI22_X1 port map( A1 => n9115, A2 => n30890, B1 => n31046, B2 => 
                           n30884, ZN => n7531);
   U24981 : OAI22_X1 port map( A1 => n9110, A2 => n30891, B1 => n31049, B2 => 
                           n30884, ZN => n7532);
   U24982 : OAI22_X1 port map( A1 => n9105, A2 => n30891, B1 => n31052, B2 => 
                           n30885, ZN => n7533);
   U24983 : OAI22_X1 port map( A1 => n9100, A2 => n30891, B1 => n31055, B2 => 
                           n30885, ZN => n7534);
   U24984 : OAI22_X1 port map( A1 => n9095, A2 => n30891, B1 => n31058, B2 => 
                           n30885, ZN => n7535);
   U24985 : OAI22_X1 port map( A1 => n9090, A2 => n30891, B1 => n31061, B2 => 
                           n30885, ZN => n7536);
   U24986 : OAI22_X1 port map( A1 => n9085, A2 => n30891, B1 => n31064, B2 => 
                           n30885, ZN => n7537);
   U24987 : OAI22_X1 port map( A1 => n9080, A2 => n30891, B1 => n31067, B2 => 
                           n30885, ZN => n7538);
   U24988 : OAI22_X1 port map( A1 => n9075, A2 => n30891, B1 => n31070, B2 => 
                           n30885, ZN => n7539);
   U24989 : OAI22_X1 port map( A1 => n9070, A2 => n30891, B1 => n31073, B2 => 
                           n30885, ZN => n7540);
   U24990 : OAI22_X1 port map( A1 => n9065, A2 => n30891, B1 => n31076, B2 => 
                           n30885, ZN => n7541);
   U24991 : OAI22_X1 port map( A1 => n9060, A2 => n30891, B1 => n31079, B2 => 
                           n30885, ZN => n7542);
   U24992 : OAI22_X1 port map( A1 => n9055, A2 => n30891, B1 => n31082, B2 => 
                           n30885, ZN => n7543);
   U24993 : OAI22_X1 port map( A1 => n9050, A2 => n30892, B1 => n31085, B2 => 
                           n30885, ZN => n7544);
   U24994 : OAI22_X1 port map( A1 => n9045, A2 => n30892, B1 => n31088, B2 => 
                           n30886, ZN => n7545);
   U24995 : OAI22_X1 port map( A1 => n9040, A2 => n30892, B1 => n31091, B2 => 
                           n30886, ZN => n7546);
   U24996 : OAI22_X1 port map( A1 => n9035, A2 => n30892, B1 => n31094, B2 => 
                           n30886, ZN => n7547);
   U24997 : OAI22_X1 port map( A1 => n9030, A2 => n30892, B1 => n31097, B2 => 
                           n30886, ZN => n7548);
   U24998 : OAI22_X1 port map( A1 => n9025, A2 => n30892, B1 => n31100, B2 => 
                           n30886, ZN => n7549);
   U24999 : OAI22_X1 port map( A1 => n9020, A2 => n30892, B1 => n31103, B2 => 
                           n30886, ZN => n7550);
   U25000 : OAI22_X1 port map( A1 => n9015, A2 => n30892, B1 => n31106, B2 => 
                           n30886, ZN => n7551);
   U25001 : OAI22_X1 port map( A1 => n9010, A2 => n30892, B1 => n31109, B2 => 
                           n30886, ZN => n7552);
   U25002 : OAI22_X1 port map( A1 => n9005, A2 => n30892, B1 => n31112, B2 => 
                           n30886, ZN => n7553);
   U25003 : OAI22_X1 port map( A1 => n9000, A2 => n30892, B1 => n31115, B2 => 
                           n30886, ZN => n7554);
   U25004 : OAI22_X1 port map( A1 => n8995, A2 => n30892, B1 => n31118, B2 => 
                           n30886, ZN => n7555);
   U25005 : OAI22_X1 port map( A1 => n8990, A2 => n30893, B1 => n31121, B2 => 
                           n30886, ZN => n7556);
   U25006 : OAI22_X1 port map( A1 => n9998, A2 => n30904, B1 => n30977, B2 => 
                           n30894, ZN => n7572);
   U25007 : OAI22_X1 port map( A1 => n9993, A2 => n30904, B1 => n30980, B2 => 
                           n30895, ZN => n7573);
   U25008 : OAI22_X1 port map( A1 => n9988, A2 => n30904, B1 => n30983, B2 => 
                           n30895, ZN => n7574);
   U25009 : OAI22_X1 port map( A1 => n9983, A2 => n30904, B1 => n30986, B2 => 
                           n30895, ZN => n7575);
   U25010 : OAI22_X1 port map( A1 => n9978, A2 => n30904, B1 => n30989, B2 => 
                           n30895, ZN => n7576);
   U25011 : OAI22_X1 port map( A1 => n9973, A2 => n30904, B1 => n30992, B2 => 
                           n30895, ZN => n7577);
   U25012 : OAI22_X1 port map( A1 => n9968, A2 => n30903, B1 => n30995, B2 => 
                           n30895, ZN => n7578);
   U25013 : OAI22_X1 port map( A1 => n9963, A2 => n30903, B1 => n30998, B2 => 
                           n30895, ZN => n7579);
   U25014 : OAI22_X1 port map( A1 => n9958, A2 => n30903, B1 => n31001, B2 => 
                           n30895, ZN => n7580);
   U25015 : OAI22_X1 port map( A1 => n9953, A2 => n30903, B1 => n31004, B2 => 
                           n30895, ZN => n7581);
   U25016 : OAI22_X1 port map( A1 => n9948, A2 => n30903, B1 => n31007, B2 => 
                           n30895, ZN => n7582);
   U25017 : OAI22_X1 port map( A1 => n9943, A2 => n30903, B1 => n31010, B2 => 
                           n30895, ZN => n7583);
   U25018 : OAI22_X1 port map( A1 => n9938, A2 => n30903, B1 => n31013, B2 => 
                           n30895, ZN => n7584);
   U25019 : OAI22_X1 port map( A1 => n9933, A2 => n30903, B1 => n31016, B2 => 
                           n30896, ZN => n7585);
   U25020 : OAI22_X1 port map( A1 => n9928, A2 => n30903, B1 => n31019, B2 => 
                           n30896, ZN => n7586);
   U25021 : OAI22_X1 port map( A1 => n9923, A2 => n30903, B1 => n31022, B2 => 
                           n30896, ZN => n7587);
   U25022 : OAI22_X1 port map( A1 => n9918, A2 => n30903, B1 => n31025, B2 => 
                           n30896, ZN => n7588);
   U25023 : OAI22_X1 port map( A1 => n9913, A2 => n30903, B1 => n31028, B2 => 
                           n30896, ZN => n7589);
   U25024 : OAI22_X1 port map( A1 => n9908, A2 => n30902, B1 => n31031, B2 => 
                           n30896, ZN => n7590);
   U25025 : OAI22_X1 port map( A1 => n9903, A2 => n30902, B1 => n31034, B2 => 
                           n30896, ZN => n7591);
   U25026 : OAI22_X1 port map( A1 => n9898, A2 => n30902, B1 => n31037, B2 => 
                           n30896, ZN => n7592);
   U25027 : OAI22_X1 port map( A1 => n9893, A2 => n30902, B1 => n31040, B2 => 
                           n30896, ZN => n7593);
   U25028 : OAI22_X1 port map( A1 => n9888, A2 => n30902, B1 => n31043, B2 => 
                           n30896, ZN => n7594);
   U25029 : OAI22_X1 port map( A1 => n9883, A2 => n30902, B1 => n31046, B2 => 
                           n30896, ZN => n7595);
   U25030 : OAI22_X1 port map( A1 => n9878, A2 => n30902, B1 => n31049, B2 => 
                           n30896, ZN => n7596);
   U25031 : OAI22_X1 port map( A1 => n9873, A2 => n30902, B1 => n31052, B2 => 
                           n30897, ZN => n7597);
   U25032 : OAI22_X1 port map( A1 => n9868, A2 => n30902, B1 => n31055, B2 => 
                           n30897, ZN => n7598);
   U25033 : OAI22_X1 port map( A1 => n9863, A2 => n30902, B1 => n31058, B2 => 
                           n30897, ZN => n7599);
   U25034 : OAI22_X1 port map( A1 => n9858, A2 => n30902, B1 => n31061, B2 => 
                           n30897, ZN => n7600);
   U25035 : OAI22_X1 port map( A1 => n9853, A2 => n30901, B1 => n31064, B2 => 
                           n30897, ZN => n7601);
   U25036 : OAI22_X1 port map( A1 => n9848, A2 => n30901, B1 => n31067, B2 => 
                           n30897, ZN => n7602);
   U25037 : OAI22_X1 port map( A1 => n9843, A2 => n30901, B1 => n31070, B2 => 
                           n30897, ZN => n7603);
   U25038 : OAI22_X1 port map( A1 => n9838, A2 => n30901, B1 => n31073, B2 => 
                           n30897, ZN => n7604);
   U25039 : OAI22_X1 port map( A1 => n9833, A2 => n30901, B1 => n31076, B2 => 
                           n30897, ZN => n7605);
   U25040 : OAI22_X1 port map( A1 => n9828, A2 => n30901, B1 => n31079, B2 => 
                           n30897, ZN => n7606);
   U25041 : OAI22_X1 port map( A1 => n9823, A2 => n30901, B1 => n31082, B2 => 
                           n30897, ZN => n7607);
   U25042 : OAI22_X1 port map( A1 => n9818, A2 => n30901, B1 => n31085, B2 => 
                           n30897, ZN => n7608);
   U25043 : OAI22_X1 port map( A1 => n9813, A2 => n30901, B1 => n31088, B2 => 
                           n30898, ZN => n7609);
   U25044 : OAI22_X1 port map( A1 => n9808, A2 => n30901, B1 => n31091, B2 => 
                           n30898, ZN => n7610);
   U25045 : OAI22_X1 port map( A1 => n9803, A2 => n30901, B1 => n31094, B2 => 
                           n30898, ZN => n7611);
   U25046 : OAI22_X1 port map( A1 => n9798, A2 => n30901, B1 => n31097, B2 => 
                           n30898, ZN => n7612);
   U25047 : OAI22_X1 port map( A1 => n9793, A2 => n30900, B1 => n31100, B2 => 
                           n30898, ZN => n7613);
   U25048 : OAI22_X1 port map( A1 => n9788, A2 => n30900, B1 => n31103, B2 => 
                           n30898, ZN => n7614);
   U25049 : OAI22_X1 port map( A1 => n9783, A2 => n30900, B1 => n31106, B2 => 
                           n30898, ZN => n7615);
   U25050 : OAI22_X1 port map( A1 => n9778, A2 => n30900, B1 => n31109, B2 => 
                           n30898, ZN => n7616);
   U25051 : OAI22_X1 port map( A1 => n9773, A2 => n30900, B1 => n31112, B2 => 
                           n30898, ZN => n7617);
   U25052 : OAI22_X1 port map( A1 => n9768, A2 => n30900, B1 => n31115, B2 => 
                           n30898, ZN => n7618);
   U25053 : OAI22_X1 port map( A1 => n9763, A2 => n30900, B1 => n31118, B2 => 
                           n30898, ZN => n7619);
   U25054 : OAI22_X1 port map( A1 => n9758, A2 => n30900, B1 => n31121, B2 => 
                           n30898, ZN => n7620);
   U25055 : OAI22_X1 port map( A1 => n30914, A2 => n25368, B1 => n30944, B2 => 
                           n30906, ZN => n7625);
   U25056 : OAI22_X1 port map( A1 => n30914, A2 => n25367, B1 => n30947, B2 => 
                           n30906, ZN => n7626);
   U25057 : OAI22_X1 port map( A1 => n30914, A2 => n25366, B1 => n30950, B2 => 
                           n30906, ZN => n7627);
   U25058 : OAI22_X1 port map( A1 => n30914, A2 => n25365, B1 => n30953, B2 => 
                           n30906, ZN => n7628);
   U25059 : OAI22_X1 port map( A1 => n30914, A2 => n25364, B1 => n30956, B2 => 
                           n30906, ZN => n7629);
   U25060 : OAI22_X1 port map( A1 => n30914, A2 => n25363, B1 => n30959, B2 => 
                           n30906, ZN => n7630);
   U25061 : OAI22_X1 port map( A1 => n30914, A2 => n25362, B1 => n30962, B2 => 
                           n30906, ZN => n7631);
   U25062 : OAI22_X1 port map( A1 => n30914, A2 => n25361, B1 => n30965, B2 => 
                           n30906, ZN => n7632);
   U25063 : OAI22_X1 port map( A1 => n30914, A2 => n25360, B1 => n30968, B2 => 
                           n30906, ZN => n7633);
   U25064 : OAI22_X1 port map( A1 => n30914, A2 => n25359, B1 => n30971, B2 => 
                           n30906, ZN => n7634);
   U25065 : OAI22_X1 port map( A1 => n30914, A2 => n25358, B1 => n30974, B2 => 
                           n30906, ZN => n7635);
   U25066 : OAI22_X1 port map( A1 => n30914, A2 => n25357, B1 => n30977, B2 => 
                           n30906, ZN => n7636);
   U25067 : OAI22_X1 port map( A1 => n30915, A2 => n25356, B1 => n30980, B2 => 
                           n30907, ZN => n7637);
   U25068 : OAI22_X1 port map( A1 => n30915, A2 => n25355, B1 => n30983, B2 => 
                           n30907, ZN => n7638);
   U25069 : OAI22_X1 port map( A1 => n30915, A2 => n25354, B1 => n30986, B2 => 
                           n30907, ZN => n7639);
   U25070 : OAI22_X1 port map( A1 => n30915, A2 => n25353, B1 => n30989, B2 => 
                           n30907, ZN => n7640);
   U25071 : OAI22_X1 port map( A1 => n30915, A2 => n25352, B1 => n30992, B2 => 
                           n30907, ZN => n7641);
   U25072 : OAI22_X1 port map( A1 => n30915, A2 => n25351, B1 => n30995, B2 => 
                           n30907, ZN => n7642);
   U25073 : OAI22_X1 port map( A1 => n30915, A2 => n25350, B1 => n30998, B2 => 
                           n30907, ZN => n7643);
   U25074 : OAI22_X1 port map( A1 => n30915, A2 => n25349, B1 => n31001, B2 => 
                           n30907, ZN => n7644);
   U25075 : OAI22_X1 port map( A1 => n30915, A2 => n25348, B1 => n31004, B2 => 
                           n30907, ZN => n7645);
   U25076 : OAI22_X1 port map( A1 => n30915, A2 => n25347, B1 => n31007, B2 => 
                           n30907, ZN => n7646);
   U25077 : OAI22_X1 port map( A1 => n30915, A2 => n25346, B1 => n31010, B2 => 
                           n30907, ZN => n7647);
   U25078 : OAI22_X1 port map( A1 => n30915, A2 => n25345, B1 => n31013, B2 => 
                           n30907, ZN => n7648);
   U25079 : OAI22_X1 port map( A1 => n30915, A2 => n25344, B1 => n31016, B2 => 
                           n30908, ZN => n7649);
   U25080 : OAI22_X1 port map( A1 => n30916, A2 => n25343, B1 => n31019, B2 => 
                           n30908, ZN => n7650);
   U25081 : OAI22_X1 port map( A1 => n30916, A2 => n25342, B1 => n31022, B2 => 
                           n30908, ZN => n7651);
   U25082 : OAI22_X1 port map( A1 => n30916, A2 => n25341, B1 => n31025, B2 => 
                           n30908, ZN => n7652);
   U25083 : OAI22_X1 port map( A1 => n30916, A2 => n25340, B1 => n31028, B2 => 
                           n30908, ZN => n7653);
   U25084 : OAI22_X1 port map( A1 => n30916, A2 => n25339, B1 => n31031, B2 => 
                           n30908, ZN => n7654);
   U25085 : OAI22_X1 port map( A1 => n30916, A2 => n25338, B1 => n31034, B2 => 
                           n30908, ZN => n7655);
   U25086 : OAI22_X1 port map( A1 => n30916, A2 => n25337, B1 => n31037, B2 => 
                           n30908, ZN => n7656);
   U25087 : OAI22_X1 port map( A1 => n30916, A2 => n25336, B1 => n31040, B2 => 
                           n30908, ZN => n7657);
   U25088 : OAI22_X1 port map( A1 => n30916, A2 => n25335, B1 => n31043, B2 => 
                           n30908, ZN => n7658);
   U25089 : OAI22_X1 port map( A1 => n30916, A2 => n25334, B1 => n31046, B2 => 
                           n30908, ZN => n7659);
   U25090 : OAI22_X1 port map( A1 => n30916, A2 => n25333, B1 => n31049, B2 => 
                           n30908, ZN => n7660);
   U25091 : OAI22_X1 port map( A1 => n30916, A2 => n25332, B1 => n31052, B2 => 
                           n30909, ZN => n7661);
   U25092 : OAI22_X1 port map( A1 => n30916, A2 => n25331, B1 => n31055, B2 => 
                           n30909, ZN => n7662);
   U25093 : OAI22_X1 port map( A1 => n30917, A2 => n25330, B1 => n31058, B2 => 
                           n30909, ZN => n7663);
   U25094 : OAI22_X1 port map( A1 => n30917, A2 => n25329, B1 => n31061, B2 => 
                           n30909, ZN => n7664);
   U25095 : OAI22_X1 port map( A1 => n30917, A2 => n25328, B1 => n31064, B2 => 
                           n30909, ZN => n7665);
   U25096 : OAI22_X1 port map( A1 => n30917, A2 => n25327, B1 => n31067, B2 => 
                           n30909, ZN => n7666);
   U25097 : OAI22_X1 port map( A1 => n30917, A2 => n25326, B1 => n31070, B2 => 
                           n30909, ZN => n7667);
   U25098 : OAI22_X1 port map( A1 => n30917, A2 => n25325, B1 => n31073, B2 => 
                           n30909, ZN => n7668);
   U25099 : OAI22_X1 port map( A1 => n30917, A2 => n25324, B1 => n31076, B2 => 
                           n30909, ZN => n7669);
   U25100 : OAI22_X1 port map( A1 => n30917, A2 => n25323, B1 => n31079, B2 => 
                           n30909, ZN => n7670);
   U25101 : OAI22_X1 port map( A1 => n30917, A2 => n25322, B1 => n31082, B2 => 
                           n30909, ZN => n7671);
   U25102 : OAI22_X1 port map( A1 => n30917, A2 => n25321, B1 => n31085, B2 => 
                           n30909, ZN => n7672);
   U25103 : OAI22_X1 port map( A1 => n30917, A2 => n25320, B1 => n31088, B2 => 
                           n30910, ZN => n7673);
   U25104 : OAI22_X1 port map( A1 => n30917, A2 => n25319, B1 => n31091, B2 => 
                           n30910, ZN => n7674);
   U25105 : OAI22_X1 port map( A1 => n30917, A2 => n25318, B1 => n31094, B2 => 
                           n30910, ZN => n7675);
   U25106 : OAI22_X1 port map( A1 => n30918, A2 => n25317, B1 => n31097, B2 => 
                           n30910, ZN => n7676);
   U25107 : OAI22_X1 port map( A1 => n30918, A2 => n25316, B1 => n31100, B2 => 
                           n30910, ZN => n7677);
   U25108 : OAI22_X1 port map( A1 => n30918, A2 => n25315, B1 => n31103, B2 => 
                           n30910, ZN => n7678);
   U25109 : OAI22_X1 port map( A1 => n30918, A2 => n25314, B1 => n31106, B2 => 
                           n30910, ZN => n7679);
   U25110 : OAI22_X1 port map( A1 => n30918, A2 => n25313, B1 => n31109, B2 => 
                           n30910, ZN => n7680);
   U25111 : OAI22_X1 port map( A1 => n30918, A2 => n25312, B1 => n31112, B2 => 
                           n30910, ZN => n7681);
   U25112 : OAI22_X1 port map( A1 => n30918, A2 => n25311, B1 => n31115, B2 => 
                           n30910, ZN => n7682);
   U25113 : OAI22_X1 port map( A1 => n30918, A2 => n25310, B1 => n31118, B2 => 
                           n30910, ZN => n7683);
   U25114 : OAI22_X1 port map( A1 => n30918, A2 => n25309, B1 => n31121, B2 => 
                           n30910, ZN => n7684);
   U25115 : OAI22_X1 port map( A1 => n9284, A2 => n30938, B1 => n30944, B2 => 
                           n30932, ZN => n7753);
   U25116 : OAI22_X1 port map( A1 => n9279, A2 => n30938, B1 => n30947, B2 => 
                           n30932, ZN => n7754);
   U25117 : OAI22_X1 port map( A1 => n9274, A2 => n30938, B1 => n30950, B2 => 
                           n30932, ZN => n7755);
   U25118 : OAI22_X1 port map( A1 => n9269, A2 => n30938, B1 => n30953, B2 => 
                           n30932, ZN => n7756);
   U25119 : OAI22_X1 port map( A1 => n9264, A2 => n30938, B1 => n30956, B2 => 
                           n30932, ZN => n7757);
   U25120 : OAI22_X1 port map( A1 => n9259, A2 => n30938, B1 => n30959, B2 => 
                           n30932, ZN => n7758);
   U25121 : OAI22_X1 port map( A1 => n9254, A2 => n30938, B1 => n30962, B2 => 
                           n30932, ZN => n7759);
   U25122 : OAI22_X1 port map( A1 => n9249, A2 => n30938, B1 => n30965, B2 => 
                           n30932, ZN => n7760);
   U25123 : OAI22_X1 port map( A1 => n9244, A2 => n30938, B1 => n30968, B2 => 
                           n30932, ZN => n7761);
   U25124 : OAI22_X1 port map( A1 => n9239, A2 => n30938, B1 => n30971, B2 => 
                           n30932, ZN => n7762);
   U25125 : OAI22_X1 port map( A1 => n9234, A2 => n30938, B1 => n30974, B2 => 
                           n30932, ZN => n7763);
   U25126 : OAI22_X1 port map( A1 => n9229, A2 => n30939, B1 => n30977, B2 => 
                           n30932, ZN => n7764);
   U25127 : OAI22_X1 port map( A1 => n9224, A2 => n30939, B1 => n30980, B2 => 
                           n30933, ZN => n7765);
   U25128 : OAI22_X1 port map( A1 => n9219, A2 => n30939, B1 => n30983, B2 => 
                           n30933, ZN => n7766);
   U25129 : OAI22_X1 port map( A1 => n9214, A2 => n30939, B1 => n30986, B2 => 
                           n30933, ZN => n7767);
   U25130 : OAI22_X1 port map( A1 => n9209, A2 => n30939, B1 => n30989, B2 => 
                           n30933, ZN => n7768);
   U25131 : OAI22_X1 port map( A1 => n9204, A2 => n30939, B1 => n30992, B2 => 
                           n30933, ZN => n7769);
   U25132 : OAI22_X1 port map( A1 => n9199, A2 => n30939, B1 => n30995, B2 => 
                           n30933, ZN => n7770);
   U25133 : OAI22_X1 port map( A1 => n9194, A2 => n30939, B1 => n30998, B2 => 
                           n30933, ZN => n7771);
   U25134 : OAI22_X1 port map( A1 => n9189, A2 => n30939, B1 => n31001, B2 => 
                           n30933, ZN => n7772);
   U25135 : OAI22_X1 port map( A1 => n9184, A2 => n30939, B1 => n31004, B2 => 
                           n30933, ZN => n7773);
   U25136 : OAI22_X1 port map( A1 => n9179, A2 => n30939, B1 => n31007, B2 => 
                           n30933, ZN => n7774);
   U25137 : OAI22_X1 port map( A1 => n9174, A2 => n30939, B1 => n31010, B2 => 
                           n30933, ZN => n7775);
   U25138 : OAI22_X1 port map( A1 => n9169, A2 => n30940, B1 => n31013, B2 => 
                           n30933, ZN => n7776);
   U25139 : OAI22_X1 port map( A1 => n9164, A2 => n30940, B1 => n31016, B2 => 
                           n30934, ZN => n7777);
   U25140 : OAI22_X1 port map( A1 => n9159, A2 => n30940, B1 => n31019, B2 => 
                           n30934, ZN => n7778);
   U25141 : OAI22_X1 port map( A1 => n9154, A2 => n30940, B1 => n31022, B2 => 
                           n30934, ZN => n7779);
   U25142 : OAI22_X1 port map( A1 => n9149, A2 => n30940, B1 => n31025, B2 => 
                           n30934, ZN => n7780);
   U25143 : OAI22_X1 port map( A1 => n9144, A2 => n30940, B1 => n31028, B2 => 
                           n30934, ZN => n7781);
   U25144 : OAI22_X1 port map( A1 => n9139, A2 => n30940, B1 => n31031, B2 => 
                           n30934, ZN => n7782);
   U25145 : OAI22_X1 port map( A1 => n9134, A2 => n30940, B1 => n31034, B2 => 
                           n30934, ZN => n7783);
   U25146 : OAI22_X1 port map( A1 => n9129, A2 => n30940, B1 => n31037, B2 => 
                           n30934, ZN => n7784);
   U25147 : OAI22_X1 port map( A1 => n9124, A2 => n30940, B1 => n31040, B2 => 
                           n30934, ZN => n7785);
   U25148 : OAI22_X1 port map( A1 => n9119, A2 => n30940, B1 => n31043, B2 => 
                           n30934, ZN => n7786);
   U25149 : OAI22_X1 port map( A1 => n9114, A2 => n30940, B1 => n31046, B2 => 
                           n30934, ZN => n7787);
   U25150 : OAI22_X1 port map( A1 => n9109, A2 => n30941, B1 => n31049, B2 => 
                           n30934, ZN => n7788);
   U25151 : OAI22_X1 port map( A1 => n9104, A2 => n30941, B1 => n31052, B2 => 
                           n30935, ZN => n7789);
   U25152 : OAI22_X1 port map( A1 => n9099, A2 => n30941, B1 => n31055, B2 => 
                           n30935, ZN => n7790);
   U25153 : OAI22_X1 port map( A1 => n9094, A2 => n30941, B1 => n31058, B2 => 
                           n30935, ZN => n7791);
   U25154 : OAI22_X1 port map( A1 => n9089, A2 => n30941, B1 => n31061, B2 => 
                           n30935, ZN => n7792);
   U25155 : OAI22_X1 port map( A1 => n9084, A2 => n30941, B1 => n31064, B2 => 
                           n30935, ZN => n7793);
   U25156 : OAI22_X1 port map( A1 => n9079, A2 => n30941, B1 => n31067, B2 => 
                           n30935, ZN => n7794);
   U25157 : OAI22_X1 port map( A1 => n9074, A2 => n30941, B1 => n31070, B2 => 
                           n30935, ZN => n7795);
   U25158 : OAI22_X1 port map( A1 => n9069, A2 => n30941, B1 => n31073, B2 => 
                           n30935, ZN => n7796);
   U25159 : OAI22_X1 port map( A1 => n9064, A2 => n30941, B1 => n31076, B2 => 
                           n30935, ZN => n7797);
   U25160 : OAI22_X1 port map( A1 => n9059, A2 => n30941, B1 => n31079, B2 => 
                           n30935, ZN => n7798);
   U25161 : OAI22_X1 port map( A1 => n9054, A2 => n30941, B1 => n31082, B2 => 
                           n30935, ZN => n7799);
   U25162 : OAI22_X1 port map( A1 => n9049, A2 => n30942, B1 => n31085, B2 => 
                           n30935, ZN => n7800);
   U25163 : OAI22_X1 port map( A1 => n9044, A2 => n30942, B1 => n31088, B2 => 
                           n30936, ZN => n7801);
   U25164 : OAI22_X1 port map( A1 => n9039, A2 => n30942, B1 => n31091, B2 => 
                           n30936, ZN => n7802);
   U25165 : OAI22_X1 port map( A1 => n9034, A2 => n30942, B1 => n31094, B2 => 
                           n30936, ZN => n7803);
   U25166 : OAI22_X1 port map( A1 => n9029, A2 => n30942, B1 => n31097, B2 => 
                           n30936, ZN => n7804);
   U25167 : OAI22_X1 port map( A1 => n9024, A2 => n30942, B1 => n31100, B2 => 
                           n30936, ZN => n7805);
   U25168 : OAI22_X1 port map( A1 => n9019, A2 => n30942, B1 => n31103, B2 => 
                           n30936, ZN => n7806);
   U25169 : OAI22_X1 port map( A1 => n9014, A2 => n30942, B1 => n31106, B2 => 
                           n30936, ZN => n7807);
   U25170 : OAI22_X1 port map( A1 => n9009, A2 => n30942, B1 => n31109, B2 => 
                           n30936, ZN => n7808);
   U25171 : OAI22_X1 port map( A1 => n9004, A2 => n30942, B1 => n31112, B2 => 
                           n30936, ZN => n7809);
   U25172 : OAI22_X1 port map( A1 => n8999, A2 => n30942, B1 => n31115, B2 => 
                           n30936, ZN => n7810);
   U25173 : OAI22_X1 port map( A1 => n8994, A2 => n30942, B1 => n31118, B2 => 
                           n30936, ZN => n7811);
   U25174 : OAI22_X1 port map( A1 => n8989, A2 => n30943, B1 => n31121, B2 => 
                           n30936, ZN => n7812);
   U25175 : OAI22_X1 port map( A1 => n9997, A2 => n31146, B1 => n31136, B2 => 
                           n30977, ZN => n7828);
   U25176 : INV_X1 port map( A => ADD_WR(1), ZN => n26101);
   U25177 : OAI221_X1 port map( B1 => n31019, B2 => n30552, C1 => n31183, C2 =>
                           n10799, A => n27341, ZN => n5819);
   U25178 : OAI21_X1 port map( B1 => n27342, B2 => n27343, A => n30546, ZN => 
                           n27341);
   U25179 : NAND4_X1 port map( A1 => n27352, A2 => n27353, A3 => n27354, A4 => 
                           n27355, ZN => n27342);
   U25180 : NAND4_X1 port map( A1 => n27344, A2 => n27345, A3 => n27346, A4 => 
                           n27347, ZN => n27343);
   U25181 : OAI221_X1 port map( B1 => n31022, B2 => n30552, C1 => n31183, C2 =>
                           n10798, A => n27315, ZN => n5821);
   U25182 : OAI21_X1 port map( B1 => n27316, B2 => n27317, A => n30546, ZN => 
                           n27315);
   U25183 : NAND4_X1 port map( A1 => n27326, A2 => n27327, A3 => n27328, A4 => 
                           n27329, ZN => n27316);
   U25184 : NAND4_X1 port map( A1 => n27318, A2 => n27319, A3 => n27320, A4 => 
                           n27321, ZN => n27317);
   U25185 : OAI221_X1 port map( B1 => n31025, B2 => n30552, C1 => n31183, C2 =>
                           n10797, A => n27289, ZN => n5823);
   U25186 : OAI21_X1 port map( B1 => n27290, B2 => n27291, A => n30546, ZN => 
                           n27289);
   U25187 : NAND4_X1 port map( A1 => n27300, A2 => n27301, A3 => n27302, A4 => 
                           n27303, ZN => n27290);
   U25188 : NAND4_X1 port map( A1 => n27292, A2 => n27293, A3 => n27294, A4 => 
                           n27295, ZN => n27291);
   U25189 : OAI221_X1 port map( B1 => n31028, B2 => n30552, C1 => n31183, C2 =>
                           n10796, A => n27263, ZN => n5825);
   U25190 : OAI21_X1 port map( B1 => n27264, B2 => n27265, A => n30546, ZN => 
                           n27263);
   U25191 : NAND4_X1 port map( A1 => n27274, A2 => n27275, A3 => n27276, A4 => 
                           n27277, ZN => n27264);
   U25192 : NAND4_X1 port map( A1 => n27266, A2 => n27267, A3 => n27268, A4 => 
                           n27269, ZN => n27265);
   U25193 : OAI221_X1 port map( B1 => n31031, B2 => n30552, C1 => n31183, C2 =>
                           n10795, A => n27237, ZN => n5827);
   U25194 : OAI21_X1 port map( B1 => n27238, B2 => n27239, A => n30546, ZN => 
                           n27237);
   U25195 : NAND4_X1 port map( A1 => n27248, A2 => n27249, A3 => n27250, A4 => 
                           n27251, ZN => n27238);
   U25196 : NAND4_X1 port map( A1 => n27240, A2 => n27241, A3 => n27242, A4 => 
                           n27243, ZN => n27239);
   U25197 : OAI221_X1 port map( B1 => n31034, B2 => n30552, C1 => n31183, C2 =>
                           n10794, A => n27211, ZN => n5829);
   U25198 : OAI21_X1 port map( B1 => n27212, B2 => n27213, A => n30546, ZN => 
                           n27211);
   U25199 : NAND4_X1 port map( A1 => n27222, A2 => n27223, A3 => n27224, A4 => 
                           n27225, ZN => n27212);
   U25200 : NAND4_X1 port map( A1 => n27214, A2 => n27215, A3 => n27216, A4 => 
                           n27217, ZN => n27213);
   U25201 : OAI221_X1 port map( B1 => n31037, B2 => n30552, C1 => n31183, C2 =>
                           n10793, A => n27185, ZN => n5831);
   U25202 : OAI21_X1 port map( B1 => n27186, B2 => n27187, A => n30546, ZN => 
                           n27185);
   U25203 : NAND4_X1 port map( A1 => n27196, A2 => n27197, A3 => n27198, A4 => 
                           n27199, ZN => n27186);
   U25204 : NAND4_X1 port map( A1 => n27188, A2 => n27189, A3 => n27190, A4 => 
                           n27191, ZN => n27187);
   U25205 : OAI221_X1 port map( B1 => n31040, B2 => n30552, C1 => n31183, C2 =>
                           n10792, A => n27159, ZN => n5833);
   U25206 : OAI21_X1 port map( B1 => n27160, B2 => n27161, A => n30546, ZN => 
                           n27159);
   U25207 : NAND4_X1 port map( A1 => n27170, A2 => n27171, A3 => n27172, A4 => 
                           n27173, ZN => n27160);
   U25208 : NAND4_X1 port map( A1 => n27162, A2 => n27163, A3 => n27164, A4 => 
                           n27165, ZN => n27161);
   U25209 : OAI221_X1 port map( B1 => n31043, B2 => n30552, C1 => n31183, C2 =>
                           n10791, A => n27133, ZN => n5835);
   U25210 : OAI21_X1 port map( B1 => n27134, B2 => n27135, A => n30546, ZN => 
                           n27133);
   U25211 : NAND4_X1 port map( A1 => n27144, A2 => n27145, A3 => n27146, A4 => 
                           n27147, ZN => n27134);
   U25212 : NAND4_X1 port map( A1 => n27136, A2 => n27137, A3 => n27138, A4 => 
                           n27139, ZN => n27135);
   U25213 : OAI221_X1 port map( B1 => n31046, B2 => n30552, C1 => n31183, C2 =>
                           n10790, A => n27107, ZN => n5837);
   U25214 : OAI21_X1 port map( B1 => n27108, B2 => n27109, A => n30546, ZN => 
                           n27107);
   U25215 : NAND4_X1 port map( A1 => n27118, A2 => n27119, A3 => n27120, A4 => 
                           n27121, ZN => n27108);
   U25216 : NAND4_X1 port map( A1 => n27110, A2 => n27111, A3 => n27112, A4 => 
                           n27113, ZN => n27109);
   U25217 : OAI221_X1 port map( B1 => n31049, B2 => n30552, C1 => n31183, C2 =>
                           n10789, A => n27081, ZN => n5839);
   U25218 : OAI21_X1 port map( B1 => n27082, B2 => n27083, A => n30546, ZN => 
                           n27081);
   U25219 : NAND4_X1 port map( A1 => n27092, A2 => n27093, A3 => n27094, A4 => 
                           n27095, ZN => n27082);
   U25220 : NAND4_X1 port map( A1 => n27084, A2 => n27085, A3 => n27086, A4 => 
                           n27087, ZN => n27083);
   U25221 : OAI221_X1 port map( B1 => n31052, B2 => n30553, C1 => n31183, C2 =>
                           n10788, A => n27055, ZN => n5841);
   U25222 : OAI21_X1 port map( B1 => n27056, B2 => n27057, A => n30547, ZN => 
                           n27055);
   U25223 : NAND4_X1 port map( A1 => n27066, A2 => n27067, A3 => n27068, A4 => 
                           n27069, ZN => n27056);
   U25224 : NAND4_X1 port map( A1 => n27058, A2 => n27059, A3 => n27060, A4 => 
                           n27061, ZN => n27057);
   U25225 : OAI221_X1 port map( B1 => n31055, B2 => n30553, C1 => n31182, C2 =>
                           n10787, A => n27029, ZN => n5843);
   U25226 : OAI21_X1 port map( B1 => n27030, B2 => n27031, A => n30547, ZN => 
                           n27029);
   U25227 : NAND4_X1 port map( A1 => n27040, A2 => n27041, A3 => n27042, A4 => 
                           n27043, ZN => n27030);
   U25228 : NAND4_X1 port map( A1 => n27032, A2 => n27033, A3 => n27034, A4 => 
                           n27035, ZN => n27031);
   U25229 : OAI221_X1 port map( B1 => n31058, B2 => n30553, C1 => n31182, C2 =>
                           n10786, A => n27003, ZN => n5845);
   U25230 : OAI21_X1 port map( B1 => n27004, B2 => n27005, A => n30547, ZN => 
                           n27003);
   U25231 : NAND4_X1 port map( A1 => n27014, A2 => n27015, A3 => n27016, A4 => 
                           n27017, ZN => n27004);
   U25232 : NAND4_X1 port map( A1 => n27006, A2 => n27007, A3 => n27008, A4 => 
                           n27009, ZN => n27005);
   U25233 : OAI221_X1 port map( B1 => n31061, B2 => n30553, C1 => n31182, C2 =>
                           n10785, A => n26977, ZN => n5847);
   U25234 : OAI21_X1 port map( B1 => n26978, B2 => n26979, A => n30547, ZN => 
                           n26977);
   U25235 : NAND4_X1 port map( A1 => n26988, A2 => n26989, A3 => n26990, A4 => 
                           n26991, ZN => n26978);
   U25236 : NAND4_X1 port map( A1 => n26980, A2 => n26981, A3 => n26982, A4 => 
                           n26983, ZN => n26979);
   U25237 : OAI221_X1 port map( B1 => n31064, B2 => n30553, C1 => n31182, C2 =>
                           n10784, A => n26951, ZN => n5849);
   U25238 : OAI21_X1 port map( B1 => n26952, B2 => n26953, A => n30547, ZN => 
                           n26951);
   U25239 : NAND4_X1 port map( A1 => n26962, A2 => n26963, A3 => n26964, A4 => 
                           n26965, ZN => n26952);
   U25240 : NAND4_X1 port map( A1 => n26954, A2 => n26955, A3 => n26956, A4 => 
                           n26957, ZN => n26953);
   U25241 : OAI221_X1 port map( B1 => n31067, B2 => n30553, C1 => n31182, C2 =>
                           n10783, A => n26925, ZN => n5851);
   U25242 : OAI21_X1 port map( B1 => n26926, B2 => n26927, A => n30547, ZN => 
                           n26925);
   U25243 : NAND4_X1 port map( A1 => n26936, A2 => n26937, A3 => n26938, A4 => 
                           n26939, ZN => n26926);
   U25244 : NAND4_X1 port map( A1 => n26928, A2 => n26929, A3 => n26930, A4 => 
                           n26931, ZN => n26927);
   U25245 : OAI221_X1 port map( B1 => n31070, B2 => n30553, C1 => n31182, C2 =>
                           n10782, A => n26899, ZN => n5853);
   U25246 : OAI21_X1 port map( B1 => n26900, B2 => n26901, A => n30547, ZN => 
                           n26899);
   U25247 : NAND4_X1 port map( A1 => n26910, A2 => n26911, A3 => n26912, A4 => 
                           n26913, ZN => n26900);
   U25248 : NAND4_X1 port map( A1 => n26902, A2 => n26903, A3 => n26904, A4 => 
                           n26905, ZN => n26901);
   U25249 : OAI221_X1 port map( B1 => n31073, B2 => n30553, C1 => n31182, C2 =>
                           n10781, A => n26873, ZN => n5855);
   U25250 : OAI21_X1 port map( B1 => n26874, B2 => n26875, A => n30547, ZN => 
                           n26873);
   U25251 : NAND4_X1 port map( A1 => n26884, A2 => n26885, A3 => n26886, A4 => 
                           n26887, ZN => n26874);
   U25252 : NAND4_X1 port map( A1 => n26876, A2 => n26877, A3 => n26878, A4 => 
                           n26879, ZN => n26875);
   U25253 : OAI221_X1 port map( B1 => n31076, B2 => n30553, C1 => n31182, C2 =>
                           n10780, A => n26847, ZN => n5857);
   U25254 : OAI21_X1 port map( B1 => n26848, B2 => n26849, A => n30547, ZN => 
                           n26847);
   U25255 : NAND4_X1 port map( A1 => n26858, A2 => n26859, A3 => n26860, A4 => 
                           n26861, ZN => n26848);
   U25256 : NAND4_X1 port map( A1 => n26850, A2 => n26851, A3 => n26852, A4 => 
                           n26853, ZN => n26849);
   U25257 : OAI221_X1 port map( B1 => n31079, B2 => n30553, C1 => n31182, C2 =>
                           n10779, A => n26821, ZN => n5859);
   U25258 : OAI21_X1 port map( B1 => n26822, B2 => n26823, A => n30547, ZN => 
                           n26821);
   U25259 : NAND4_X1 port map( A1 => n26832, A2 => n26833, A3 => n26834, A4 => 
                           n26835, ZN => n26822);
   U25260 : NAND4_X1 port map( A1 => n26824, A2 => n26825, A3 => n26826, A4 => 
                           n26827, ZN => n26823);
   U25261 : OAI221_X1 port map( B1 => n31082, B2 => n30553, C1 => n31182, C2 =>
                           n10778, A => n26795, ZN => n5861);
   U25262 : OAI21_X1 port map( B1 => n26796, B2 => n26797, A => n30547, ZN => 
                           n26795);
   U25263 : NAND4_X1 port map( A1 => n26806, A2 => n26807, A3 => n26808, A4 => 
                           n26809, ZN => n26796);
   U25264 : NAND4_X1 port map( A1 => n26798, A2 => n26799, A3 => n26800, A4 => 
                           n26801, ZN => n26797);
   U25265 : OAI221_X1 port map( B1 => n31085, B2 => n30553, C1 => n31182, C2 =>
                           n10777, A => n26769, ZN => n5863);
   U25266 : OAI21_X1 port map( B1 => n26770, B2 => n26771, A => n30547, ZN => 
                           n26769);
   U25267 : NAND4_X1 port map( A1 => n26780, A2 => n26781, A3 => n26782, A4 => 
                           n26783, ZN => n26770);
   U25268 : NAND4_X1 port map( A1 => n26772, A2 => n26773, A3 => n26774, A4 => 
                           n26775, ZN => n26771);
   U25269 : OAI221_X1 port map( B1 => n31088, B2 => n30554, C1 => n31182, C2 =>
                           n10776, A => n26743, ZN => n5865);
   U25270 : OAI21_X1 port map( B1 => n26744, B2 => n26745, A => n30548, ZN => 
                           n26743);
   U25271 : NAND4_X1 port map( A1 => n26754, A2 => n26755, A3 => n26756, A4 => 
                           n26757, ZN => n26744);
   U25272 : NAND4_X1 port map( A1 => n26746, A2 => n26747, A3 => n26748, A4 => 
                           n26749, ZN => n26745);
   U25273 : OAI221_X1 port map( B1 => n31091, B2 => n30554, C1 => n31182, C2 =>
                           n10775, A => n26717, ZN => n5867);
   U25274 : OAI21_X1 port map( B1 => n26718, B2 => n26719, A => n30548, ZN => 
                           n26717);
   U25275 : NAND4_X1 port map( A1 => n26728, A2 => n26729, A3 => n26730, A4 => 
                           n26731, ZN => n26718);
   U25276 : NAND4_X1 port map( A1 => n26720, A2 => n26721, A3 => n26722, A4 => 
                           n26723, ZN => n26719);
   U25277 : OAI221_X1 port map( B1 => n31094, B2 => n30554, C1 => n31181, C2 =>
                           n10774, A => n26691, ZN => n5869);
   U25278 : OAI21_X1 port map( B1 => n26692, B2 => n26693, A => n30548, ZN => 
                           n26691);
   U25279 : NAND4_X1 port map( A1 => n26702, A2 => n26703, A3 => n26704, A4 => 
                           n26705, ZN => n26692);
   U25280 : NAND4_X1 port map( A1 => n26694, A2 => n26695, A3 => n26696, A4 => 
                           n26697, ZN => n26693);
   U25281 : OAI221_X1 port map( B1 => n31097, B2 => n30554, C1 => n31181, C2 =>
                           n10773, A => n26665, ZN => n5871);
   U25282 : OAI21_X1 port map( B1 => n26666, B2 => n26667, A => n30548, ZN => 
                           n26665);
   U25283 : NAND4_X1 port map( A1 => n26676, A2 => n26677, A3 => n26678, A4 => 
                           n26679, ZN => n26666);
   U25284 : NAND4_X1 port map( A1 => n26668, A2 => n26669, A3 => n26670, A4 => 
                           n26671, ZN => n26667);
   U25285 : OAI221_X1 port map( B1 => n31100, B2 => n30554, C1 => n31181, C2 =>
                           n10772, A => n26639, ZN => n5873);
   U25286 : OAI21_X1 port map( B1 => n26640, B2 => n26641, A => n30548, ZN => 
                           n26639);
   U25287 : NAND4_X1 port map( A1 => n26650, A2 => n26651, A3 => n26652, A4 => 
                           n26653, ZN => n26640);
   U25288 : NAND4_X1 port map( A1 => n26642, A2 => n26643, A3 => n26644, A4 => 
                           n26645, ZN => n26641);
   U25289 : OAI221_X1 port map( B1 => n31103, B2 => n30554, C1 => n31181, C2 =>
                           n10771, A => n26613, ZN => n5875);
   U25290 : OAI21_X1 port map( B1 => n26614, B2 => n26615, A => n30548, ZN => 
                           n26613);
   U25291 : NAND4_X1 port map( A1 => n26624, A2 => n26625, A3 => n26626, A4 => 
                           n26627, ZN => n26614);
   U25292 : NAND4_X1 port map( A1 => n26616, A2 => n26617, A3 => n26618, A4 => 
                           n26619, ZN => n26615);
   U25293 : OAI221_X1 port map( B1 => n31106, B2 => n30554, C1 => n31181, C2 =>
                           n10770, A => n26587, ZN => n5877);
   U25294 : OAI21_X1 port map( B1 => n26588, B2 => n26589, A => n30548, ZN => 
                           n26587);
   U25295 : NAND4_X1 port map( A1 => n26598, A2 => n26599, A3 => n26600, A4 => 
                           n26601, ZN => n26588);
   U25296 : NAND4_X1 port map( A1 => n26590, A2 => n26591, A3 => n26592, A4 => 
                           n26593, ZN => n26589);
   U25297 : OAI221_X1 port map( B1 => n31109, B2 => n30554, C1 => n31181, C2 =>
                           n10769, A => n26561, ZN => n5879);
   U25298 : OAI21_X1 port map( B1 => n26562, B2 => n26563, A => n30548, ZN => 
                           n26561);
   U25299 : NAND4_X1 port map( A1 => n26572, A2 => n26573, A3 => n26574, A4 => 
                           n26575, ZN => n26562);
   U25300 : NAND4_X1 port map( A1 => n26564, A2 => n26565, A3 => n26566, A4 => 
                           n26567, ZN => n26563);
   U25301 : OAI221_X1 port map( B1 => n31112, B2 => n30554, C1 => n31181, C2 =>
                           n10768, A => n26535, ZN => n5881);
   U25302 : OAI21_X1 port map( B1 => n26536, B2 => n26537, A => n30548, ZN => 
                           n26535);
   U25303 : NAND4_X1 port map( A1 => n26546, A2 => n26547, A3 => n26548, A4 => 
                           n26549, ZN => n26536);
   U25304 : NAND4_X1 port map( A1 => n26538, A2 => n26539, A3 => n26540, A4 => 
                           n26541, ZN => n26537);
   U25305 : OAI221_X1 port map( B1 => n31115, B2 => n30554, C1 => n31181, C2 =>
                           n10767, A => n26509, ZN => n5883);
   U25306 : OAI21_X1 port map( B1 => n26510, B2 => n26511, A => n30548, ZN => 
                           n26509);
   U25307 : NAND4_X1 port map( A1 => n26520, A2 => n26521, A3 => n26522, A4 => 
                           n26523, ZN => n26510);
   U25308 : NAND4_X1 port map( A1 => n26512, A2 => n26513, A3 => n26514, A4 => 
                           n26515, ZN => n26511);
   U25309 : OAI221_X1 port map( B1 => n31118, B2 => n30554, C1 => n31181, C2 =>
                           n10766, A => n26483, ZN => n5885);
   U25310 : OAI21_X1 port map( B1 => n26484, B2 => n26485, A => n30548, ZN => 
                           n26483);
   U25311 : NAND4_X1 port map( A1 => n26494, A2 => n26495, A3 => n26496, A4 => 
                           n26497, ZN => n26484);
   U25312 : NAND4_X1 port map( A1 => n26486, A2 => n26487, A3 => n26488, A4 => 
                           n26489, ZN => n26485);
   U25313 : OAI221_X1 port map( B1 => n31121, B2 => n30554, C1 => n31181, C2 =>
                           n10765, A => n26457, ZN => n5887);
   U25314 : OAI21_X1 port map( B1 => n26458, B2 => n26459, A => n30548, ZN => 
                           n26457);
   U25315 : NAND4_X1 port map( A1 => n26468, A2 => n26469, A3 => n26470, A4 => 
                           n26471, ZN => n26458);
   U25316 : NAND4_X1 port map( A1 => n26460, A2 => n26461, A3 => n26462, A4 => 
                           n26463, ZN => n26459);
   U25317 : INV_X1 port map( A => ADD_RD1(3), ZN => n29293);
   U25318 : INV_X1 port map( A => ADD_RD2(0), ZN => n28007);
   U25319 : OAI221_X1 port map( B1 => n31124, B2 => n30350, C1 => n31185, C2 =>
                           n10828, A => n28132, ZN => n5762);
   U25320 : OAI21_X1 port map( B1 => n28133, B2 => n28134, A => n30344, ZN => 
                           n28132);
   U25321 : NAND4_X1 port map( A1 => n28135, A2 => n28136, A3 => n28137, A4 => 
                           n28138, ZN => n28134);
   U25322 : NAND4_X1 port map( A1 => n28143, A2 => n28144, A3 => n28145, A4 => 
                           n28146, ZN => n28133);
   U25323 : OAI221_X1 port map( B1 => n31127, B2 => n30350, C1 => n31186, C2 =>
                           n10827, A => n28113, ZN => n5764);
   U25324 : OAI21_X1 port map( B1 => n28114, B2 => n28115, A => n30344, ZN => 
                           n28113);
   U25325 : NAND4_X1 port map( A1 => n28116, A2 => n28117, A3 => n28118, A4 => 
                           n28119, ZN => n28115);
   U25326 : NAND4_X1 port map( A1 => n28124, A2 => n28125, A3 => n28126, A4 => 
                           n28127, ZN => n28114);
   U25327 : OAI221_X1 port map( B1 => n31130, B2 => n30350, C1 => n31185, C2 =>
                           n10826, A => n28094, ZN => n5766);
   U25328 : OAI21_X1 port map( B1 => n28095, B2 => n28096, A => n30344, ZN => 
                           n28094);
   U25329 : NAND4_X1 port map( A1 => n28097, A2 => n28098, A3 => n28099, A4 => 
                           n28100, ZN => n28096);
   U25330 : NAND4_X1 port map( A1 => n28105, A2 => n28106, A3 => n28107, A4 => 
                           n28108, ZN => n28095);
   U25331 : OAI221_X1 port map( B1 => n31133, B2 => n30350, C1 => n31186, C2 =>
                           n10825, A => n28041, ZN => n5768);
   U25332 : OAI21_X1 port map( B1 => n28042, B2 => n28043, A => n30344, ZN => 
                           n28041);
   U25333 : NAND4_X1 port map( A1 => n28045, A2 => n28046, A3 => n28047, A4 => 
                           n28048, ZN => n28043);
   U25334 : NAND4_X1 port map( A1 => n28069, A2 => n28070, A3 => n28071, A4 => 
                           n28072, ZN => n28042);
   U25335 : OAI221_X1 port map( B1 => n30944, B2 => n30550, C1 => n31185, C2 =>
                           n10824, A => n27991, ZN => n5769);
   U25336 : OAI21_X1 port map( B1 => n27992, B2 => n27993, A => n30544, ZN => 
                           n27991);
   U25337 : NAND4_X1 port map( A1 => n27995, A2 => n27996, A3 => n27997, A4 => 
                           n27998, ZN => n27993);
   U25338 : NAND4_X1 port map( A1 => n28014, A2 => n28015, A3 => n28016, A4 => 
                           n28017, ZN => n27992);
   U25339 : OAI221_X1 port map( B1 => n30947, B2 => n30550, C1 => n31185, C2 =>
                           n10823, A => n27965, ZN => n5771);
   U25340 : OAI21_X1 port map( B1 => n27966, B2 => n27967, A => n30544, ZN => 
                           n27965);
   U25341 : NAND4_X1 port map( A1 => n27968, A2 => n27969, A3 => n27970, A4 => 
                           n27971, ZN => n27967);
   U25342 : NAND4_X1 port map( A1 => n27976, A2 => n27977, A3 => n27978, A4 => 
                           n27979, ZN => n27966);
   U25343 : OAI221_X1 port map( B1 => n30950, B2 => n30550, C1 => n31185, C2 =>
                           n10822, A => n27939, ZN => n5773);
   U25344 : OAI21_X1 port map( B1 => n27940, B2 => n27941, A => n30544, ZN => 
                           n27939);
   U25345 : NAND4_X1 port map( A1 => n27942, A2 => n27943, A3 => n27944, A4 => 
                           n27945, ZN => n27941);
   U25346 : NAND4_X1 port map( A1 => n27950, A2 => n27951, A3 => n27952, A4 => 
                           n27953, ZN => n27940);
   U25347 : OAI221_X1 port map( B1 => n30953, B2 => n30550, C1 => n31185, C2 =>
                           n10821, A => n27913, ZN => n5775);
   U25348 : OAI21_X1 port map( B1 => n27914, B2 => n27915, A => n30544, ZN => 
                           n27913);
   U25349 : NAND4_X1 port map( A1 => n27916, A2 => n27917, A3 => n27918, A4 => 
                           n27919, ZN => n27915);
   U25350 : NAND4_X1 port map( A1 => n27924, A2 => n27925, A3 => n27926, A4 => 
                           n27927, ZN => n27914);
   U25351 : OAI221_X1 port map( B1 => n30956, B2 => n30550, C1 => n31185, C2 =>
                           n10820, A => n27887, ZN => n5777);
   U25352 : OAI21_X1 port map( B1 => n27888, B2 => n27889, A => n30544, ZN => 
                           n27887);
   U25353 : NAND4_X1 port map( A1 => n27890, A2 => n27891, A3 => n27892, A4 => 
                           n27893, ZN => n27889);
   U25354 : NAND4_X1 port map( A1 => n27898, A2 => n27899, A3 => n27900, A4 => 
                           n27901, ZN => n27888);
   U25355 : OAI221_X1 port map( B1 => n30959, B2 => n30550, C1 => n31185, C2 =>
                           n10819, A => n27861, ZN => n5779);
   U25356 : OAI21_X1 port map( B1 => n27862, B2 => n27863, A => n30544, ZN => 
                           n27861);
   U25357 : NAND4_X1 port map( A1 => n27864, A2 => n27865, A3 => n27866, A4 => 
                           n27867, ZN => n27863);
   U25358 : NAND4_X1 port map( A1 => n27872, A2 => n27873, A3 => n27874, A4 => 
                           n27875, ZN => n27862);
   U25359 : OAI221_X1 port map( B1 => n30962, B2 => n30550, C1 => n31185, C2 =>
                           n10818, A => n27835, ZN => n5781);
   U25360 : OAI21_X1 port map( B1 => n27836, B2 => n27837, A => n30544, ZN => 
                           n27835);
   U25361 : NAND4_X1 port map( A1 => n27838, A2 => n27839, A3 => n27840, A4 => 
                           n27841, ZN => n27837);
   U25362 : NAND4_X1 port map( A1 => n27846, A2 => n27847, A3 => n27848, A4 => 
                           n27849, ZN => n27836);
   U25363 : OAI221_X1 port map( B1 => n30965, B2 => n30550, C1 => n31185, C2 =>
                           n10817, A => n27809, ZN => n5783);
   U25364 : OAI21_X1 port map( B1 => n27810, B2 => n27811, A => n30544, ZN => 
                           n27809);
   U25365 : NAND4_X1 port map( A1 => n27812, A2 => n27813, A3 => n27814, A4 => 
                           n27815, ZN => n27811);
   U25366 : NAND4_X1 port map( A1 => n27820, A2 => n27821, A3 => n27822, A4 => 
                           n27823, ZN => n27810);
   U25367 : OAI221_X1 port map( B1 => n30968, B2 => n30550, C1 => n31185, C2 =>
                           n10816, A => n27783, ZN => n5785);
   U25368 : OAI21_X1 port map( B1 => n27784, B2 => n27785, A => n30544, ZN => 
                           n27783);
   U25369 : NAND4_X1 port map( A1 => n27786, A2 => n27787, A3 => n27788, A4 => 
                           n27789, ZN => n27785);
   U25370 : NAND4_X1 port map( A1 => n27794, A2 => n27795, A3 => n27796, A4 => 
                           n27797, ZN => n27784);
   U25371 : OAI221_X1 port map( B1 => n30971, B2 => n30550, C1 => n31185, C2 =>
                           n10815, A => n27757, ZN => n5787);
   U25372 : OAI21_X1 port map( B1 => n27758, B2 => n27759, A => n30544, ZN => 
                           n27757);
   U25373 : NAND4_X1 port map( A1 => n27760, A2 => n27761, A3 => n27762, A4 => 
                           n27763, ZN => n27759);
   U25374 : NAND4_X1 port map( A1 => n27768, A2 => n27769, A3 => n27770, A4 => 
                           n27771, ZN => n27758);
   U25375 : OAI221_X1 port map( B1 => n30974, B2 => n30550, C1 => n31185, C2 =>
                           n10814, A => n27731, ZN => n5789);
   U25376 : OAI21_X1 port map( B1 => n27732, B2 => n27733, A => n30544, ZN => 
                           n27731);
   U25377 : NAND4_X1 port map( A1 => n27734, A2 => n27735, A3 => n27736, A4 => 
                           n27737, ZN => n27733);
   U25378 : NAND4_X1 port map( A1 => n27742, A2 => n27743, A3 => n27744, A4 => 
                           n27745, ZN => n27732);
   U25379 : OAI221_X1 port map( B1 => n30977, B2 => n30550, C1 => n31184, C2 =>
                           n10813, A => n27705, ZN => n5791);
   U25380 : OAI21_X1 port map( B1 => n27706, B2 => n27707, A => n30544, ZN => 
                           n27705);
   U25381 : NAND4_X1 port map( A1 => n27708, A2 => n27709, A3 => n27710, A4 => 
                           n27711, ZN => n27707);
   U25382 : NAND4_X1 port map( A1 => n27716, A2 => n27717, A3 => n27718, A4 => 
                           n27719, ZN => n27706);
   U25383 : OAI221_X1 port map( B1 => n30980, B2 => n30551, C1 => n31184, C2 =>
                           n10812, A => n27679, ZN => n5793);
   U25384 : OAI21_X1 port map( B1 => n27680, B2 => n27681, A => n30545, ZN => 
                           n27679);
   U25385 : NAND4_X1 port map( A1 => n27682, A2 => n27683, A3 => n27684, A4 => 
                           n27685, ZN => n27681);
   U25386 : NAND4_X1 port map( A1 => n27690, A2 => n27691, A3 => n27692, A4 => 
                           n27693, ZN => n27680);
   U25387 : OAI221_X1 port map( B1 => n30983, B2 => n30551, C1 => n31184, C2 =>
                           n10811, A => n27653, ZN => n5795);
   U25388 : OAI21_X1 port map( B1 => n27654, B2 => n27655, A => n30545, ZN => 
                           n27653);
   U25389 : NAND4_X1 port map( A1 => n27656, A2 => n27657, A3 => n27658, A4 => 
                           n27659, ZN => n27655);
   U25390 : NAND4_X1 port map( A1 => n27664, A2 => n27665, A3 => n27666, A4 => 
                           n27667, ZN => n27654);
   U25391 : OAI221_X1 port map( B1 => n30986, B2 => n30551, C1 => n31184, C2 =>
                           n10810, A => n27627, ZN => n5797);
   U25392 : OAI21_X1 port map( B1 => n27628, B2 => n27629, A => n30545, ZN => 
                           n27627);
   U25393 : NAND4_X1 port map( A1 => n27630, A2 => n27631, A3 => n27632, A4 => 
                           n27633, ZN => n27629);
   U25394 : NAND4_X1 port map( A1 => n27638, A2 => n27639, A3 => n27640, A4 => 
                           n27641, ZN => n27628);
   U25395 : OAI221_X1 port map( B1 => n30989, B2 => n30551, C1 => n31184, C2 =>
                           n10809, A => n27601, ZN => n5799);
   U25396 : OAI21_X1 port map( B1 => n27602, B2 => n27603, A => n30545, ZN => 
                           n27601);
   U25397 : NAND4_X1 port map( A1 => n27604, A2 => n27605, A3 => n27606, A4 => 
                           n27607, ZN => n27603);
   U25398 : NAND4_X1 port map( A1 => n27612, A2 => n27613, A3 => n27614, A4 => 
                           n27615, ZN => n27602);
   U25399 : OAI221_X1 port map( B1 => n30992, B2 => n30551, C1 => n31184, C2 =>
                           n10808, A => n27575, ZN => n5801);
   U25400 : OAI21_X1 port map( B1 => n27576, B2 => n27577, A => n30545, ZN => 
                           n27575);
   U25401 : NAND4_X1 port map( A1 => n27578, A2 => n27579, A3 => n27580, A4 => 
                           n27581, ZN => n27577);
   U25402 : NAND4_X1 port map( A1 => n27586, A2 => n27587, A3 => n27588, A4 => 
                           n27589, ZN => n27576);
   U25403 : OAI221_X1 port map( B1 => n30995, B2 => n30551, C1 => n31184, C2 =>
                           n10807, A => n27549, ZN => n5803);
   U25404 : OAI21_X1 port map( B1 => n27550, B2 => n27551, A => n30545, ZN => 
                           n27549);
   U25405 : NAND4_X1 port map( A1 => n27552, A2 => n27553, A3 => n27554, A4 => 
                           n27555, ZN => n27551);
   U25406 : NAND4_X1 port map( A1 => n27560, A2 => n27561, A3 => n27562, A4 => 
                           n27563, ZN => n27550);
   U25407 : OAI221_X1 port map( B1 => n30998, B2 => n30551, C1 => n31184, C2 =>
                           n10806, A => n27523, ZN => n5805);
   U25408 : OAI21_X1 port map( B1 => n27524, B2 => n27525, A => n30545, ZN => 
                           n27523);
   U25409 : NAND4_X1 port map( A1 => n27526, A2 => n27527, A3 => n27528, A4 => 
                           n27529, ZN => n27525);
   U25410 : NAND4_X1 port map( A1 => n27534, A2 => n27535, A3 => n27536, A4 => 
                           n27537, ZN => n27524);
   U25411 : OAI221_X1 port map( B1 => n31001, B2 => n30551, C1 => n31184, C2 =>
                           n10805, A => n27497, ZN => n5807);
   U25412 : OAI21_X1 port map( B1 => n27498, B2 => n27499, A => n30545, ZN => 
                           n27497);
   U25413 : NAND4_X1 port map( A1 => n27500, A2 => n27501, A3 => n27502, A4 => 
                           n27503, ZN => n27499);
   U25414 : NAND4_X1 port map( A1 => n27508, A2 => n27509, A3 => n27510, A4 => 
                           n27511, ZN => n27498);
   U25415 : OAI221_X1 port map( B1 => n31004, B2 => n30551, C1 => n31184, C2 =>
                           n10804, A => n27471, ZN => n5809);
   U25416 : OAI21_X1 port map( B1 => n27472, B2 => n27473, A => n30545, ZN => 
                           n27471);
   U25417 : NAND4_X1 port map( A1 => n27474, A2 => n27475, A3 => n27476, A4 => 
                           n27477, ZN => n27473);
   U25418 : NAND4_X1 port map( A1 => n27482, A2 => n27483, A3 => n27484, A4 => 
                           n27485, ZN => n27472);
   U25419 : OAI221_X1 port map( B1 => n31007, B2 => n30551, C1 => n31184, C2 =>
                           n10803, A => n27445, ZN => n5811);
   U25420 : OAI21_X1 port map( B1 => n27446, B2 => n27447, A => n30545, ZN => 
                           n27445);
   U25421 : NAND4_X1 port map( A1 => n27448, A2 => n27449, A3 => n27450, A4 => 
                           n27451, ZN => n27447);
   U25422 : NAND4_X1 port map( A1 => n27456, A2 => n27457, A3 => n27458, A4 => 
                           n27459, ZN => n27446);
   U25423 : OAI221_X1 port map( B1 => n31010, B2 => n30551, C1 => n31184, C2 =>
                           n10802, A => n27419, ZN => n5813);
   U25424 : OAI21_X1 port map( B1 => n27420, B2 => n27421, A => n30545, ZN => 
                           n27419);
   U25425 : NAND4_X1 port map( A1 => n27422, A2 => n27423, A3 => n27424, A4 => 
                           n27425, ZN => n27421);
   U25426 : NAND4_X1 port map( A1 => n27430, A2 => n27431, A3 => n27432, A4 => 
                           n27433, ZN => n27420);
   U25427 : OAI221_X1 port map( B1 => n31013, B2 => n30551, C1 => n31184, C2 =>
                           n10801, A => n27393, ZN => n5815);
   U25428 : OAI21_X1 port map( B1 => n27394, B2 => n27395, A => n30545, ZN => 
                           n27393);
   U25429 : NAND4_X1 port map( A1 => n27396, A2 => n27397, A3 => n27398, A4 => 
                           n27399, ZN => n27395);
   U25430 : NAND4_X1 port map( A1 => n27404, A2 => n27405, A3 => n27406, A4 => 
                           n27407, ZN => n27394);
   U25431 : OAI221_X1 port map( B1 => n31016, B2 => n30552, C1 => n31183, C2 =>
                           n10800, A => n27367, ZN => n5817);
   U25432 : OAI21_X1 port map( B1 => n27368, B2 => n27369, A => n30546, ZN => 
                           n27367);
   U25433 : NAND4_X1 port map( A1 => n27370, A2 => n27371, A3 => n27372, A4 => 
                           n27373, ZN => n27369);
   U25434 : NAND4_X1 port map( A1 => n27378, A2 => n27379, A3 => n27380, A4 => 
                           n27381, ZN => n27368);
   U25435 : OAI221_X1 port map( B1 => n31133, B2 => n30555, C1 => n31180, C2 =>
                           n10761, A => n26320, ZN => n5895);
   U25436 : OAI21_X1 port map( B1 => n26321, B2 => n26322, A => n30549, ZN => 
                           n26320);
   U25437 : NAND4_X1 port map( A1 => n26348, A2 => n26349, A3 => n26350, A4 => 
                           n26351, ZN => n26321);
   U25438 : NAND4_X1 port map( A1 => n26324, A2 => n26325, A3 => n26326, A4 => 
                           n26327, ZN => n26322);
   U25439 : INV_X1 port map( A => ADD_RD1(0), ZN => n29288);
   U25440 : INV_X1 port map( A => ADD_RD2(3), ZN => n28024);
   U25441 : NAND4_X1 port map( A1 => n29309, A2 => n29310, A3 => n29311, A4 => 
                           n29312, ZN => n29275);
   U25442 : XNOR2_X1 port map( A => ADD_RD1(3), B => ADD_WR(3), ZN => n29309);
   U25443 : XNOR2_X1 port map( A => ADD_RD1(2), B => ADD_WR(2), ZN => n29311);
   U25444 : XNOR2_X1 port map( A => ADD_RD1(0), B => ADD_WR(0), ZN => n29310);
   U25445 : NAND4_X1 port map( A1 => n28034, A2 => n28035, A3 => n28036, A4 => 
                           n28037, ZN => n27994);
   U25446 : XNOR2_X1 port map( A => ADD_RD2(0), B => ADD_WR(0), ZN => n28034);
   U25447 : XNOR2_X1 port map( A => ADD_RD2(2), B => ADD_WR(2), ZN => n28036);
   U25448 : XNOR2_X1 port map( A => ADD_RD2(3), B => ADD_WR(3), ZN => n28035);
   U25449 : OR2_X1 port map( A1 => n29275, A2 => RESET, ZN => n28040);
   U25450 : OR2_X1 port map( A1 => n27994, A2 => RESET, ZN => n26319);
   U25451 : OAI21_X1 port map( B1 => n31174, B2 => n10980, A => n30144, ZN => 
                           n5713);
   U25452 : OAI21_X1 port map( B1 => n31174, B2 => n10979, A => n30144, ZN => 
                           n5715);
   U25453 : OAI21_X1 port map( B1 => n31171, B2 => n10978, A => n30144, ZN => 
                           n5717);
   U25454 : OAI21_X1 port map( B1 => n31170, B2 => n10977, A => n30144, ZN => 
                           n5719);
   U25455 : OAI21_X1 port map( B1 => n31170, B2 => n10976, A => n30144, ZN => 
                           n5721);
   U25456 : OAI21_X1 port map( B1 => n31170, B2 => n10975, A => n30144, ZN => 
                           n5723);
   U25457 : OAI21_X1 port map( B1 => n31171, B2 => n10974, A => n30144, ZN => 
                           n5725);
   U25458 : OAI21_X1 port map( B1 => n31172, B2 => n10973, A => n30144, ZN => 
                           n5727);
   U25459 : OAI21_X1 port map( B1 => n31173, B2 => n10972, A => n30144, ZN => 
                           n5729);
   U25460 : OAI21_X1 port map( B1 => n31173, B2 => n10971, A => n30144, ZN => 
                           n5731);
   U25461 : OAI21_X1 port map( B1 => n31174, B2 => n10970, A => n30144, ZN => 
                           n5733);
   U25462 : OAI21_X1 port map( B1 => n31174, B2 => n10969, A => n30144, ZN => 
                           n5735);
   U25463 : OAI21_X1 port map( B1 => n31171, B2 => n10968, A => n30145, ZN => 
                           n5737);
   U25464 : OAI21_X1 port map( B1 => n31171, B2 => n10967, A => n30145, ZN => 
                           n5739);
   U25465 : OAI21_X1 port map( B1 => n31171, B2 => n10966, A => n30145, ZN => 
                           n5741);
   U25466 : OAI21_X1 port map( B1 => n31170, B2 => n10965, A => n30145, ZN => 
                           n5743);
   U25467 : OAI21_X1 port map( B1 => n31170, B2 => n10964, A => n30145, ZN => 
                           n5745);
   U25468 : OAI21_X1 port map( B1 => n31170, B2 => n10963, A => n30145, ZN => 
                           n5747);
   U25469 : OAI21_X1 port map( B1 => n31167, B2 => n10962, A => n30145, ZN => 
                           n5749);
   U25470 : OAI21_X1 port map( B1 => n31163, B2 => n10961, A => n30145, ZN => 
                           n5751);
   U25471 : OAI21_X1 port map( B1 => n31164, B2 => n10960, A => n30145, ZN => 
                           n5753);
   U25472 : OAI21_X1 port map( B1 => n31163, B2 => n10959, A => n30145, ZN => 
                           n5755);
   U25473 : OAI21_X1 port map( B1 => n31164, B2 => n10958, A => n30145, ZN => 
                           n5757);
   U25474 : OAI21_X1 port map( B1 => n31164, B2 => n10957, A => n30145, ZN => 
                           n5759);
   U25475 : OAI21_X1 port map( B1 => n31167, B2 => n10916, A => n31151, ZN => 
                           n7917);
   U25476 : OAI21_X1 port map( B1 => n31167, B2 => n10915, A => n31151, ZN => 
                           n7918);
   U25477 : OAI21_X1 port map( B1 => n31165, B2 => n10914, A => n31151, ZN => 
                           n7919);
   U25478 : OAI21_X1 port map( B1 => n31168, B2 => n10913, A => n31151, ZN => 
                           n7920);
   U25479 : OAI21_X1 port map( B1 => n31168, B2 => n10912, A => n31151, ZN => 
                           n7921);
   U25480 : OAI21_X1 port map( B1 => n31168, B2 => n10911, A => n31151, ZN => 
                           n7922);
   U25481 : OAI21_X1 port map( B1 => n31168, B2 => n10910, A => n31151, ZN => 
                           n7923);
   U25482 : OAI21_X1 port map( B1 => n31168, B2 => n10909, A => n31151, ZN => 
                           n7924);
   U25483 : OAI21_X1 port map( B1 => n31168, B2 => n10908, A => n31151, ZN => 
                           n7925);
   U25484 : OAI21_X1 port map( B1 => n31168, B2 => n10907, A => n31151, ZN => 
                           n7926);
   U25485 : OAI21_X1 port map( B1 => n31168, B2 => n10906, A => n31151, ZN => 
                           n7927);
   U25486 : OAI21_X1 port map( B1 => n31168, B2 => n10905, A => n31151, ZN => 
                           n7928);
   U25487 : OAI21_X1 port map( B1 => n31168, B2 => n10904, A => n31152, ZN => 
                           n7929);
   U25488 : OAI21_X1 port map( B1 => n31168, B2 => n10903, A => n31152, ZN => 
                           n7930);
   U25489 : OAI21_X1 port map( B1 => n31168, B2 => n10902, A => n31152, ZN => 
                           n7931);
   U25490 : OAI21_X1 port map( B1 => n31169, B2 => n10901, A => n31152, ZN => 
                           n7932);
   U25491 : OAI21_X1 port map( B1 => n31169, B2 => n10900, A => n31152, ZN => 
                           n7933);
   U25492 : OAI21_X1 port map( B1 => n31169, B2 => n10899, A => n31152, ZN => 
                           n7934);
   U25493 : OAI21_X1 port map( B1 => n31169, B2 => n10898, A => n31152, ZN => 
                           n7935);
   U25494 : OAI21_X1 port map( B1 => n31169, B2 => n10897, A => n31152, ZN => 
                           n7936);
   U25495 : OAI21_X1 port map( B1 => n31169, B2 => n10896, A => n31152, ZN => 
                           n7937);
   U25496 : OAI21_X1 port map( B1 => n31169, B2 => n10895, A => n31152, ZN => 
                           n7938);
   U25497 : OAI21_X1 port map( B1 => n31169, B2 => n10894, A => n31152, ZN => 
                           n7939);
   U25498 : OAI21_X1 port map( B1 => n31169, B2 => n10893, A => n31152, ZN => 
                           n7940);
   U25499 : OAI21_X1 port map( B1 => n31164, B2 => n10956, A => n30146, ZN => 
                           n5761);
   U25500 : OAI21_X1 port map( B1 => n31164, B2 => n10955, A => n30146, ZN => 
                           n5763);
   U25501 : OAI21_X1 port map( B1 => n31164, B2 => n10954, A => n30146, ZN => 
                           n5765);
   U25502 : OAI21_X1 port map( B1 => n31164, B2 => n10953, A => n30146, ZN => 
                           n5767);
   U25503 : OAI21_X1 port map( B1 => n31169, B2 => n10892, A => n31153, ZN => 
                           n7941);
   U25504 : OAI21_X1 port map( B1 => n31169, B2 => n10891, A => n31153, ZN => 
                           n7942);
   U25505 : OAI21_X1 port map( B1 => n31169, B2 => n10890, A => n31153, ZN => 
                           n7943);
   U25506 : OAI21_X1 port map( B1 => n31170, B2 => n10889, A => n31153, ZN => 
                           n7944);
   U25507 : INV_X1 port map( A => WR, ZN => n25806);
   U25508 : AND3_X1 port map( A1 => WR, A2 => ENABLE, A3 => ADD_WR(4), ZN => 
                           n26091);
   U25509 : INV_X1 port map( A => ENABLE, ZN => n25152);
   U25510 : OAI21_X1 port map( B1 => n31164, B2 => n11016, A => n30141, ZN => 
                           n5641);
   U25511 : OAI21_X1 port map( B1 => n31170, B2 => n11015, A => n30141, ZN => 
                           n5643);
   U25512 : OAI21_X1 port map( B1 => n31170, B2 => n11014, A => n30141, ZN => 
                           n5645);
   U25513 : OAI21_X1 port map( B1 => n31170, B2 => n11013, A => n30141, ZN => 
                           n5647);
   U25514 : OAI21_X1 port map( B1 => n31171, B2 => n11012, A => n30141, ZN => 
                           n5649);
   U25515 : OAI21_X1 port map( B1 => n31170, B2 => n11011, A => n30141, ZN => 
                           n5651);
   U25516 : OAI21_X1 port map( B1 => n31170, B2 => n11010, A => n30141, ZN => 
                           n5653);
   U25517 : OAI21_X1 port map( B1 => n31171, B2 => n11009, A => n30141, ZN => 
                           n5655);
   U25518 : OAI21_X1 port map( B1 => n31171, B2 => n11008, A => n30141, ZN => 
                           n5657);
   U25519 : OAI21_X1 port map( B1 => n31172, B2 => n11007, A => n30141, ZN => 
                           n5659);
   U25520 : OAI21_X1 port map( B1 => n31172, B2 => n11006, A => n30141, ZN => 
                           n5661);
   U25521 : OAI21_X1 port map( B1 => n31172, B2 => n11005, A => n30141, ZN => 
                           n5663);
   U25522 : OAI21_X1 port map( B1 => n31172, B2 => n11004, A => n30142, ZN => 
                           n5665);
   U25523 : OAI21_X1 port map( B1 => n31172, B2 => n11003, A => n30142, ZN => 
                           n5667);
   U25524 : OAI21_X1 port map( B1 => n31171, B2 => n11002, A => n30142, ZN => 
                           n5669);
   U25525 : OAI21_X1 port map( B1 => n31171, B2 => n11001, A => n30142, ZN => 
                           n5671);
   U25526 : OAI21_X1 port map( B1 => n31172, B2 => n11000, A => n30142, ZN => 
                           n5673);
   U25527 : OAI21_X1 port map( B1 => n31172, B2 => n10999, A => n30142, ZN => 
                           n5675);
   U25528 : OAI21_X1 port map( B1 => n31171, B2 => n10998, A => n30142, ZN => 
                           n5677);
   U25529 : OAI21_X1 port map( B1 => n31172, B2 => n10997, A => n30142, ZN => 
                           n5679);
   U25530 : OAI21_X1 port map( B1 => n31172, B2 => n10996, A => n30142, ZN => 
                           n5681);
   U25531 : OAI21_X1 port map( B1 => n31171, B2 => n10995, A => n30142, ZN => 
                           n5683);
   U25532 : OAI21_X1 port map( B1 => n31173, B2 => n10994, A => n30142, ZN => 
                           n5685);
   U25533 : OAI21_X1 port map( B1 => n31173, B2 => n10993, A => n30142, ZN => 
                           n5687);
   U25534 : OAI21_X1 port map( B1 => n31172, B2 => n10992, A => n30143, ZN => 
                           n5689);
   U25535 : OAI21_X1 port map( B1 => n31173, B2 => n10991, A => n30143, ZN => 
                           n5691);
   U25536 : OAI21_X1 port map( B1 => n31173, B2 => n10990, A => n30143, ZN => 
                           n5693);
   U25537 : OAI21_X1 port map( B1 => n31172, B2 => n10989, A => n30143, ZN => 
                           n5695);
   U25538 : OAI21_X1 port map( B1 => n31173, B2 => n10988, A => n30143, ZN => 
                           n5697);
   U25539 : OAI21_X1 port map( B1 => n31173, B2 => n10987, A => n30143, ZN => 
                           n5699);
   U25540 : OAI21_X1 port map( B1 => n31173, B2 => n10986, A => n30143, ZN => 
                           n5701);
   U25541 : OAI21_X1 port map( B1 => n31173, B2 => n10985, A => n30143, ZN => 
                           n5703);
   U25542 : OAI21_X1 port map( B1 => n31173, B2 => n10984, A => n30143, ZN => 
                           n5705);
   U25543 : OAI21_X1 port map( B1 => n31173, B2 => n10982, A => n30143, ZN => 
                           n5709);
   U25544 : OAI21_X1 port map( B1 => n31164, B2 => n10952, A => n31148, ZN => 
                           n7881);
   U25545 : OAI21_X1 port map( B1 => n31164, B2 => n10951, A => n31148, ZN => 
                           n7882);
   U25546 : OAI21_X1 port map( B1 => n31164, B2 => n10950, A => n31148, ZN => 
                           n7883);
   U25547 : OAI21_X1 port map( B1 => n31164, B2 => n10949, A => n31148, ZN => 
                           n7884);
   U25548 : OAI21_X1 port map( B1 => n31165, B2 => n10948, A => n31148, ZN => 
                           n7885);
   U25549 : OAI21_X1 port map( B1 => n31165, B2 => n10947, A => n31148, ZN => 
                           n7886);
   U25550 : OAI21_X1 port map( B1 => n31165, B2 => n10946, A => n31148, ZN => 
                           n7887);
   U25551 : OAI21_X1 port map( B1 => n31165, B2 => n10945, A => n31148, ZN => 
                           n7888);
   U25552 : OAI21_X1 port map( B1 => n31165, B2 => n10944, A => n31148, ZN => 
                           n7889);
   U25553 : OAI21_X1 port map( B1 => n31165, B2 => n10943, A => n31148, ZN => 
                           n7890);
   U25554 : OAI21_X1 port map( B1 => n31165, B2 => n10942, A => n31148, ZN => 
                           n7891);
   U25555 : OAI21_X1 port map( B1 => n31165, B2 => n10941, A => n31148, ZN => 
                           n7892);
   U25556 : OAI21_X1 port map( B1 => n31165, B2 => n10940, A => n31149, ZN => 
                           n7893);
   U25557 : OAI21_X1 port map( B1 => n31165, B2 => n10939, A => n31149, ZN => 
                           n7894);
   U25558 : OAI21_X1 port map( B1 => n31165, B2 => n10938, A => n31149, ZN => 
                           n7895);
   U25559 : OAI21_X1 port map( B1 => n31166, B2 => n10937, A => n31149, ZN => 
                           n7896);
   U25560 : OAI21_X1 port map( B1 => n31166, B2 => n10936, A => n31149, ZN => 
                           n7897);
   U25561 : OAI21_X1 port map( B1 => n31166, B2 => n10935, A => n31149, ZN => 
                           n7898);
   U25562 : OAI21_X1 port map( B1 => n31166, B2 => n10934, A => n31149, ZN => 
                           n7899);
   U25563 : OAI21_X1 port map( B1 => n31166, B2 => n10933, A => n31149, ZN => 
                           n7900);
   U25564 : OAI21_X1 port map( B1 => n31166, B2 => n10932, A => n31149, ZN => 
                           n7901);
   U25565 : OAI21_X1 port map( B1 => n31166, B2 => n10931, A => n31149, ZN => 
                           n7902);
   U25566 : OAI21_X1 port map( B1 => n31166, B2 => n10930, A => n31149, ZN => 
                           n7903);
   U25567 : OAI21_X1 port map( B1 => n31166, B2 => n10929, A => n31149, ZN => 
                           n7904);
   U25568 : OAI21_X1 port map( B1 => n31166, B2 => n10928, A => n31150, ZN => 
                           n7905);
   U25569 : OAI21_X1 port map( B1 => n31166, B2 => n10927, A => n31150, ZN => 
                           n7906);
   U25570 : OAI21_X1 port map( B1 => n31166, B2 => n10926, A => n31150, ZN => 
                           n7907);
   U25571 : OAI21_X1 port map( B1 => n31167, B2 => n10925, A => n31150, ZN => 
                           n7908);
   U25572 : OAI21_X1 port map( B1 => n31167, B2 => n10924, A => n31150, ZN => 
                           n7909);
   U25573 : OAI21_X1 port map( B1 => n31167, B2 => n10923, A => n31150, ZN => 
                           n7910);
   U25574 : OAI21_X1 port map( B1 => n31167, B2 => n10922, A => n31150, ZN => 
                           n7911);
   U25575 : OAI21_X1 port map( B1 => n31167, B2 => n10921, A => n31150, ZN => 
                           n7912);
   U25576 : OAI21_X1 port map( B1 => n31167, B2 => n10920, A => n31150, ZN => 
                           n7913);
   U25577 : OAI21_X1 port map( B1 => n31167, B2 => n10919, A => n31150, ZN => 
                           n7914);
   U25578 : OAI21_X1 port map( B1 => n31167, B2 => n10918, A => n31150, ZN => 
                           n7915);
   U25579 : OAI21_X1 port map( B1 => n31167, B2 => n10917, A => n31150, ZN => 
                           n7916);
   U25580 : OAI21_X1 port map( B1 => n31174, B2 => n10983, A => n30143, ZN => 
                           n5707);
   U25581 : OAI21_X1 port map( B1 => n31174, B2 => n10981, A => n30143, ZN => 
                           n5711);
   U25582 : INV_X1 port map( A => DATAIN(0), ZN => n25230);
   U25583 : INV_X1 port map( A => DATAIN(1), ZN => n25228);
   U25584 : INV_X1 port map( A => DATAIN(2), ZN => n25226);
   U25585 : INV_X1 port map( A => DATAIN(3), ZN => n25224);
   U25586 : INV_X1 port map( A => DATAIN(4), ZN => n25222);
   U25587 : INV_X1 port map( A => DATAIN(5), ZN => n25220);
   U25588 : INV_X1 port map( A => DATAIN(6), ZN => n25218);
   U25589 : INV_X1 port map( A => DATAIN(7), ZN => n25216);
   U25590 : INV_X1 port map( A => DATAIN(8), ZN => n25214);
   U25591 : INV_X1 port map( A => DATAIN(9), ZN => n25212);
   U25592 : INV_X1 port map( A => DATAIN(10), ZN => n25210);
   U25593 : INV_X1 port map( A => DATAIN(11), ZN => n25208);
   U25594 : INV_X1 port map( A => DATAIN(12), ZN => n25207);
   U25595 : INV_X1 port map( A => DATAIN(13), ZN => n25206);
   U25596 : INV_X1 port map( A => DATAIN(14), ZN => n25205);
   U25597 : INV_X1 port map( A => DATAIN(15), ZN => n25204);
   U25598 : INV_X1 port map( A => DATAIN(16), ZN => n25203);
   U25599 : INV_X1 port map( A => DATAIN(17), ZN => n25202);
   U25600 : INV_X1 port map( A => DATAIN(18), ZN => n25201);
   U25601 : INV_X1 port map( A => DATAIN(19), ZN => n25200);
   U25602 : INV_X1 port map( A => DATAIN(20), ZN => n25199);
   U25603 : INV_X1 port map( A => DATAIN(21), ZN => n25198);
   U25604 : INV_X1 port map( A => DATAIN(22), ZN => n25197);
   U25605 : INV_X1 port map( A => DATAIN(23), ZN => n25196);
   U25606 : INV_X1 port map( A => DATAIN(24), ZN => n25195);
   U25607 : INV_X1 port map( A => DATAIN(25), ZN => n25194);
   U25608 : INV_X1 port map( A => DATAIN(26), ZN => n25193);
   U25609 : INV_X1 port map( A => DATAIN(27), ZN => n25192);
   U25610 : INV_X1 port map( A => DATAIN(28), ZN => n25191);
   U25611 : INV_X1 port map( A => DATAIN(29), ZN => n25190);
   U25612 : INV_X1 port map( A => DATAIN(30), ZN => n25189);
   U25613 : INV_X1 port map( A => DATAIN(31), ZN => n25188);
   U25614 : INV_X1 port map( A => DATAIN(32), ZN => n25187);
   U25615 : INV_X1 port map( A => DATAIN(33), ZN => n25186);
   U25616 : INV_X1 port map( A => DATAIN(34), ZN => n25185);
   U25617 : INV_X1 port map( A => DATAIN(35), ZN => n25184);
   U25618 : INV_X1 port map( A => DATAIN(36), ZN => n25183);
   U25619 : INV_X1 port map( A => DATAIN(37), ZN => n25182);
   U25620 : INV_X1 port map( A => DATAIN(38), ZN => n25181);
   U25621 : INV_X1 port map( A => DATAIN(39), ZN => n25180);
   U25622 : INV_X1 port map( A => DATAIN(40), ZN => n25179);
   U25623 : INV_X1 port map( A => DATAIN(41), ZN => n25178);
   U25624 : INV_X1 port map( A => DATAIN(42), ZN => n25177);
   U25625 : INV_X1 port map( A => DATAIN(43), ZN => n25176);
   U25626 : INV_X1 port map( A => DATAIN(44), ZN => n25175);
   U25627 : INV_X1 port map( A => DATAIN(45), ZN => n25174);
   U25628 : INV_X1 port map( A => DATAIN(46), ZN => n25173);
   U25629 : INV_X1 port map( A => DATAIN(47), ZN => n25172);
   U25630 : INV_X1 port map( A => DATAIN(48), ZN => n25171);
   U25631 : INV_X1 port map( A => DATAIN(49), ZN => n25170);
   U25632 : INV_X1 port map( A => DATAIN(50), ZN => n25169);
   U25633 : INV_X1 port map( A => DATAIN(51), ZN => n25168);
   U25634 : INV_X1 port map( A => DATAIN(52), ZN => n25167);
   U25635 : INV_X1 port map( A => DATAIN(53), ZN => n25166);
   U25636 : INV_X1 port map( A => DATAIN(54), ZN => n25165);
   U25637 : INV_X1 port map( A => DATAIN(55), ZN => n25164);
   U25638 : INV_X1 port map( A => DATAIN(56), ZN => n25163);
   U25639 : INV_X1 port map( A => DATAIN(57), ZN => n25162);
   U25640 : INV_X1 port map( A => DATAIN(58), ZN => n25161);
   U25641 : INV_X1 port map( A => DATAIN(59), ZN => n25160);
   U25642 : INV_X1 port map( A => DATAIN(60), ZN => n25159);
   U25643 : INV_X1 port map( A => DATAIN(61), ZN => n25158);
   U25644 : INV_X1 port map( A => DATAIN(62), ZN => n25157);
   U25645 : INV_X1 port map( A => DATAIN(63), ZN => n25156);
   U25646 : INV_X1 port map( A => ADD_WR(3), ZN => n25453);
   U25647 : INV_X1 port map( A => ADD_WR(0), ZN => n25452);
   U25648 : INV_X1 port map( A => RD1, ZN => n29313);
   U25649 : INV_X1 port map( A => RD2, ZN => n25153);
   U25650 : INV_X1 port map( A => ADD_RD1(1), ZN => n29308);
   U25651 : INV_X1 port map( A => ADD_RD2(1), ZN => n28033);
   U25652 : INV_X1 port map( A => ADD_RD1(2), ZN => n29305);
   U25653 : INV_X1 port map( A => ADD_RD2(2), ZN => n28028);
   U25654 : INV_X1 port map( A => ADD_WR(2), ZN => n26100);
   U25655 : INV_X1 port map( A => RESET, ZN => n25150);
   U25656 : CLKBUF_X1 port map( A => n28093, Z => n30146);
   U25657 : CLKBUF_X1 port map( A => n28092, Z => n30152);
   U25658 : CLKBUF_X1 port map( A => n28091, Z => n30158);
   U25659 : CLKBUF_X1 port map( A => n28089, Z => n30164);
   U25660 : CLKBUF_X1 port map( A => n28088, Z => n30170);
   U25661 : CLKBUF_X1 port map( A => n28087, Z => n30176);
   U25662 : CLKBUF_X1 port map( A => n28086, Z => n30182);
   U25663 : CLKBUF_X1 port map( A => n28084, Z => n30188);
   U25664 : CLKBUF_X1 port map( A => n28083, Z => n30194);
   U25665 : CLKBUF_X1 port map( A => n28082, Z => n30200);
   U25666 : CLKBUF_X1 port map( A => n28081, Z => n30206);
   U25667 : CLKBUF_X1 port map( A => n28079, Z => n30212);
   U25668 : CLKBUF_X1 port map( A => n28078, Z => n30218);
   U25669 : CLKBUF_X1 port map( A => n28077, Z => n30224);
   U25670 : CLKBUF_X1 port map( A => n28076, Z => n30230);
   U25671 : CLKBUF_X1 port map( A => n28074, Z => n30236);
   U25672 : CLKBUF_X1 port map( A => n28073, Z => n30242);
   U25673 : CLKBUF_X1 port map( A => n28068, Z => n30248);
   U25674 : CLKBUF_X1 port map( A => n28067, Z => n30254);
   U25675 : CLKBUF_X1 port map( A => n28065, Z => n30260);
   U25676 : CLKBUF_X1 port map( A => n28064, Z => n30266);
   U25677 : CLKBUF_X1 port map( A => n28063, Z => n30272);
   U25678 : CLKBUF_X1 port map( A => n28062, Z => n30278);
   U25679 : CLKBUF_X1 port map( A => n28060, Z => n30284);
   U25680 : CLKBUF_X1 port map( A => n28059, Z => n30290);
   U25681 : CLKBUF_X1 port map( A => n28058, Z => n30296);
   U25682 : CLKBUF_X1 port map( A => n28057, Z => n30302);
   U25683 : CLKBUF_X1 port map( A => n28055, Z => n30308);
   U25684 : CLKBUF_X1 port map( A => n28054, Z => n30314);
   U25685 : CLKBUF_X1 port map( A => n28053, Z => n30320);
   U25686 : CLKBUF_X1 port map( A => n28052, Z => n30326);
   U25687 : CLKBUF_X1 port map( A => n28050, Z => n30332);
   U25688 : CLKBUF_X1 port map( A => n28049, Z => n30338);
   U25689 : CLKBUF_X1 port map( A => n28044, Z => n30344);
   U25690 : CLKBUF_X1 port map( A => n28040, Z => n30350);
   U25691 : CLKBUF_X1 port map( A => n26377, Z => n30356);
   U25692 : CLKBUF_X1 port map( A => n26376, Z => n30362);
   U25693 : CLKBUF_X1 port map( A => n26373, Z => n30368);
   U25694 : CLKBUF_X1 port map( A => n26371, Z => n30374);
   U25695 : CLKBUF_X1 port map( A => n26370, Z => n30380);
   U25696 : CLKBUF_X1 port map( A => n26369, Z => n30386);
   U25697 : CLKBUF_X1 port map( A => n26366, Z => n30392);
   U25698 : CLKBUF_X1 port map( A => n26364, Z => n30398);
   U25699 : CLKBUF_X1 port map( A => n26363, Z => n30404);
   U25700 : CLKBUF_X1 port map( A => n26362, Z => n30410);
   U25701 : CLKBUF_X1 port map( A => n26359, Z => n30416);
   U25702 : CLKBUF_X1 port map( A => n26357, Z => n30422);
   U25703 : CLKBUF_X1 port map( A => n26356, Z => n30428);
   U25704 : CLKBUF_X1 port map( A => n26355, Z => n30434);
   U25705 : CLKBUF_X1 port map( A => n26353, Z => n30440);
   U25706 : CLKBUF_X1 port map( A => n26352, Z => n30446);
   U25707 : CLKBUF_X1 port map( A => n26347, Z => n30452);
   U25708 : CLKBUF_X1 port map( A => n26344, Z => n30465);
   U25709 : CLKBUF_X1 port map( A => n26343, Z => n30471);
   U25710 : CLKBUF_X1 port map( A => n26342, Z => n30477);
   U25711 : CLKBUF_X1 port map( A => n26341, Z => n30483);
   U25712 : CLKBUF_X1 port map( A => n26339, Z => n30489);
   U25713 : CLKBUF_X1 port map( A => n26338, Z => n30495);
   U25714 : CLKBUF_X1 port map( A => n26337, Z => n30501);
   U25715 : CLKBUF_X1 port map( A => n26336, Z => n30507);
   U25716 : CLKBUF_X1 port map( A => n26334, Z => n30513);
   U25717 : CLKBUF_X1 port map( A => n26333, Z => n30519);
   U25718 : CLKBUF_X1 port map( A => n26332, Z => n30525);
   U25719 : CLKBUF_X1 port map( A => n26331, Z => n30531);
   U25720 : CLKBUF_X1 port map( A => n26329, Z => n30537);
   U25721 : CLKBUF_X1 port map( A => n26328, Z => n30543);
   U25722 : CLKBUF_X1 port map( A => n26323, Z => n30549);
   U25723 : CLKBUF_X1 port map( A => n26319, Z => n30555);
   U25724 : CLKBUF_X1 port map( A => n26318, Z => n30561);
   U25725 : CLKBUF_X1 port map( A => n26252, Z => n30574);
   U25726 : CLKBUF_X1 port map( A => n26249, Z => n30587);
   U25727 : CLKBUF_X1 port map( A => n26248, Z => n30593);
   U25728 : CLKBUF_X1 port map( A => n26235, Z => n30599);
   U25729 : CLKBUF_X1 port map( A => n26234, Z => n30605);
   U25730 : CLKBUF_X1 port map( A => n26170, Z => n30611);
   U25731 : CLKBUF_X1 port map( A => n26104, Z => n30624);
   U25732 : CLKBUF_X1 port map( A => n26098, Z => n30637);
   U25733 : CLKBUF_X1 port map( A => n26097, Z => n30643);
   U25734 : CLKBUF_X1 port map( A => n26095, Z => n30649);
   U25735 : CLKBUF_X1 port map( A => n26094, Z => n30655);
   U25736 : CLKBUF_X1 port map( A => n26093, Z => n30661);
   U25737 : CLKBUF_X1 port map( A => n26092, Z => n30667);
   U25738 : CLKBUF_X1 port map( A => n26090, Z => n30673);
   U25739 : CLKBUF_X1 port map( A => n26089, Z => n30679);
   U25740 : CLKBUF_X1 port map( A => n26025, Z => n30685);
   U25741 : CLKBUF_X1 port map( A => n25959, Z => n30698);
   U25742 : CLKBUF_X1 port map( A => n25956, Z => n30711);
   U25743 : CLKBUF_X1 port map( A => n25955, Z => n30717);
   U25744 : CLKBUF_X1 port map( A => n25942, Z => n30723);
   U25745 : CLKBUF_X1 port map( A => n25941, Z => n30729);
   U25746 : CLKBUF_X1 port map( A => n25876, Z => n30735);
   U25747 : CLKBUF_X1 port map( A => n25809, Z => n30748);
   U25748 : CLKBUF_X1 port map( A => n25805, Z => n30761);
   U25749 : CLKBUF_X1 port map( A => n25804, Z => n30767);
   U25750 : CLKBUF_X1 port map( A => n25803, Z => n30773);
   U25751 : CLKBUF_X1 port map( A => n25802, Z => n30779);
   U25752 : CLKBUF_X1 port map( A => n25738, Z => n30785);
   U25753 : CLKBUF_X1 port map( A => n25672, Z => n30798);
   U25754 : CLKBUF_X1 port map( A => n25669, Z => n30811);
   U25755 : CLKBUF_X1 port map( A => n25668, Z => n30817);
   U25756 : CLKBUF_X1 port map( A => n25656, Z => n30823);
   U25757 : CLKBUF_X1 port map( A => n25655, Z => n30829);
   U25758 : CLKBUF_X1 port map( A => n25590, Z => n30835);
   U25759 : CLKBUF_X1 port map( A => n25523, Z => n30848);
   U25760 : CLKBUF_X1 port map( A => n25457, Z => n30861);
   U25761 : CLKBUF_X1 port map( A => n25387, Z => n30874);
   U25762 : CLKBUF_X1 port map( A => n25384, Z => n30887);
   U25763 : CLKBUF_X1 port map( A => n25383, Z => n30893);
   U25764 : CLKBUF_X1 port map( A => n25370, Z => n30899);
   U25765 : CLKBUF_X1 port map( A => n25369, Z => n30905);
   U25766 : CLKBUF_X1 port map( A => n25305, Z => n30911);
   U25767 : CLKBUF_X1 port map( A => n25238, Z => n30924);
   U25768 : CLKBUF_X1 port map( A => n25234, Z => n30937);
   U25769 : CLKBUF_X1 port map( A => n25233, Z => n30943);
   U25770 : CLKBUF_X1 port map( A => n25155, Z => n31141);
   U25771 : CLKBUF_X1 port map( A => n25154, Z => n31147);
   U25772 : CLKBUF_X1 port map( A => n25151, Z => n31153);
   U25773 : CLKBUF_X1 port map( A => n31158, Z => n31187);

end SYN_A;
